{
"addr/interpolation":[
"Adressinterpolering"
],
"address":[
"postadress",
"postnummer",
"husnummer",
"Adress",
"destination",
"gatuadress",
"adress",
"postort"
],
"advertising/billboard":[
"annonstavla",
"affischtavla",
"reklamskylt",
"reklamtavla",
"affisch",
"reklam",
"Annonstavla"
],
"advertising/board":[
"anslagstavla",
"tillkännagivanden",
"Anslagstavla",
"reklam",
"reklamblad",
"korktavla",
"whiteboard",
"flygblad"
],
"advertising/column":[
"annonstavla",
"reklamplats",
"Reklampelare",
"annons",
"affisch",
"reklam",
"affischpelare",
"reklampelare",
"billboard",
"marknadsföring",
"annonspelare",
"annonsering"
],
"advertising/poster_box":[
"affischtavla",
"reklamyta",
"reklamtavla",
"reklamlåda",
"reklambox",
"reklampelare",
"Reklamtavla"
],
"advertising/totem":[
"skyltpylon",
"Skyltpylon",
"skylttavla på stolpe",
"reklam på stolpe",
"reklampelare",
"stolpskylt"
],
"aerialway":[
"Linbaneobjekt"
],
"aerialway/cable_car":[
"Kabinbana",
"linbana",
"kabinbana",
"pendelbana"
],
"aerialway/chair_lift":[
"stollift",
"expresslift",
"lift",
"linbana",
"Stollift",
"stolslift",
"skidlift"
],
"aerialway/drag_lift":[
"Släplift",
"släplift",
"lift",
"linbana",
"skidlift",
"draglift"
],
"aerialway/gondola":[
"gondol",
"lift",
"linbana",
"skidlift",
"gondolbana",
"Gondollinbana"
],
"aerialway/goods":[
"gruvlift",
"transportbana",
"varor",
"gods",
"varulift",
"linbana",
"transport",
"industrilift",
"transportlift",
"transportlinbana",
"lift",
"industri",
"Transportlinbana"
],
"aerialway/j-bar":[
"j-lift",
"ankarlift",
"j-bygellift",
"släplift",
"lift",
"linbana",
"skidlift",
"J-krokslift"
],
"aerialway/magic_carpet":[
"rullband",
"skidliften",
"släplift",
"lift",
"Rullband",
"magisk matta"
],
"aerialway/mixed_lift":[
"Hybridlift (Telemixlift)",
"stollift",
"expresslift",
"gondol",
"lift",
"linbana",
"telemixlift",
"skidlift",
"stolslift",
"hybridlift",
"gondolbana"
],
"aerialway/platter":[
"tallrikslift",
"släplift",
"lift",
"knapp",
"knapplift",
"linbana",
"tallrik",
"skidlift",
"Knapplift"
],
"aerialway/pylon":[
"pylon",
"stolpe",
"Linbanestolpe",
"stötta",
"pelare"
],
"aerialway/rope_tow":[
"replift",
"släplift",
"lift",
"linbana",
"skidlift",
"Replift"
],
"aerialway/t-bar":[
"Ankarlift",
"ankarlift",
"t-bygellift",
"släplift",
"lift",
"t-lift",
"linbana",
"skidlift"
],
"aerialway/zip_line":[
"zipwire",
"glidbana",
"zipline",
"zip-line",
"linbana",
"travers",
"Zipline"
],
"aeroway":[
"Flygtrafiksobjekt"
],
"aeroway/aerodrome":[
"flyghamn",
"flyg",
"flygplats",
"aerodrom",
"Flygplats",
"lufthamn",
"flygfält",
"flygplan",
"landningsplats"
],
"aeroway/apron":[
"Parkering för flygplan (Apron)",
"tamac",
"ramp",
"flygparkering",
"parkering av flygplan",
"apron",
"parkering av plan",
"flygplansplatta",
"flygplatsplatta",
"flygplansparkering",
"taxibana"
],
"aeroway/gate":[
"flyggate",
"flygplatsgate",
"Gate",
"gate"
],
"aeroway/hangar":[
"hangar",
"flygverkstad",
"Hangar",
"flygplansgarage",
"flyggarage",
"garage för flygplan",
"flygplanshall"
],
"aeroway/helipad":[
"helikopterplatta",
"Helikopterplatta",
"helikopter",
"helipad"
],
"aeroway/holding_position":[
"holding",
"ils",
"väntplats",
"väntplats för flygplan",
"holding position",
"mls",
"Väntplats för flygplan"
],
"aeroway/jet_bridge":[
"jetbridge",
"landgång",
"pbb",
"brygga",
"Ombordstigningsbrygga",
"passagerarbrygga",
"skybridge",
"jet bridge",
"gate",
"ombordstigningsbrygga",
"embarkeringsbrygga"
],
"aeroway/parking_position":[
"flyg",
"flygparkering",
"flygplan",
"parkeringsplats för flygplan",
"parkering",
"Parkeringsplats för flygplan"
],
"aeroway/runway":[
"Start- och landningsbana",
"flyg",
"rwy",
"flygplats",
"landningsbana",
"landa",
"landning",
"landningsfällt",
"startbana",
"rullbana"
],
"aeroway/spaceport":[
"raketuppsättningssida",
"rymdport",
"avfyrningsplats. raketramp",
"raketuppskjutningscenter",
"raketuppskattningskomplex",
"raketuppskjutning",
"kosmodrom",
"rymdbas",
"raketområde",
"Rymdbas",
"raket"
],
"aeroway/taxiway":[
"flygplansväg",
"transportbana",
"taxiway",
"transportsträcka",
"Taxibana",
"taxibana"
],
"aeroway/terminal":[
"flygplats",
"Flygterminal",
"flygterminal",
"terminal",
"avgångshall",
"ankomsthall",
"flygplatsterminal"
],
"aeroway/windsock":[
"Vindstrut",
"vindstrut",
"vindriktning",
"strut",
"vindmätning",
"vindstyrka",
"vind"
],
"allotments/plot":[
"odlingslott",
"lott",
"koloniträdgård",
"kolonilott",
"koloniområde",
"koloni",
"Kolonilott",
"täppa"
],
"amenity":[
"Facilitet"
],
"amenity/animal_boarding":[
"kattpensionat",
"katt",
"hundkollo",
"Djurhotell",
"katthotell",
"hundhotell",
"häst",
"hundpensionat",
"hund",
"inackordering",
"reptil",
"djurkollo",
"djurpensionat",
"djurhotell",
"husdjur",
"kattkollo"
],
"amenity/animal_breeding":[
"katt",
"ko",
"tjur",
"kattunge",
"djurhållning",
"uppfödning",
"häst",
"avel",
"hund",
"reptil",
"valp",
"boskap",
"Djuruppfödning",
"djuravel",
"husdjur",
"djuruppfödning"
],
"amenity/animal_shelter":[
"Djurhem",
"katthem",
"hemlös",
"katt",
"rovfågel",
"häst",
"vanvårdad",
"hund",
"reptil",
"omplacering",
"djuradoption",
"karantän",
"djurhem",
"husdjur",
"omhändertagande",
"djurskydd"
],
"amenity/arts_centre":[
"kulturcenter",
"konstcenter",
"museum",
"kultur",
"tavlor",
"kulturhus",
"konst",
"Konstcenter"
],
"amenity/atm":[
"bankomat",
"minuten",
"otto",
"uttagsautomat",
"Uttagsautomat",
"atm",
"kontanter",
"pengar"
],
"amenity/bank":[
"kreditinrättning",
"investering",
"Bank",
"bankkontor",
"insättning",
"check",
"låneinstitut",
"bankvalv",
"besparing",
"bank",
"penninginrättning",
"fonder",
"banklokal",
"kassa",
"penninganstalt"
],
"amenity/bar":[
"bar",
"Bar",
"matställe",
"servering",
"saloon",
"öl",
"cocktailsalong",
"sprit",
"pub",
"krog"
],
"amenity/bar/lgbtq":[
"hbtq-bar",
"lgbtq bar",
"gay-bar",
"lgb bar",
"lesbisk bar",
"lgbt bar",
"HBTQ-bar"
],
"amenity/bbq":[
"bbq",
"barbecue",
"eldning",
"eldstad",
"grillplats",
"Grillplats/Grill",
"grill",
"eldplats",
"grillning"
],
"amenity/bench":[
"sits",
"bänk",
"sittmöbel",
"sittbräde",
"soffa",
"Bänk"
],
"amenity/bicycle_parking":[
"cykelparkering",
"ställplats",
"cykel",
"Cykelparkering",
"cykelställ",
"parkering"
],
"amenity/bicycle_parking/building":[
"Cykelparkeringsgarage",
"cykelparkeringsgarage",
"cykelparkering",
"cykel",
"flervåningscykelgarage",
"garage",
"parkering",
"flervåningscykelparkering"
],
"amenity/bicycle_parking/lockers":[
"cykellås",
"fastlåsning av cykel",
"cykel",
"Cykellås",
"fastlåsning",
"lås"
],
"amenity/bicycle_parking/shed":[
"cykelskydd",
"cykelparkering",
"cykelparkeringsskydd",
"Cykelskydd",
"cykel",
"cykeltak",
"tak",
"cykelparkeringstak"
],
"amenity/bicycle_rental":[
"Cykeluthyrning",
"lånecykel",
"cykellån",
"cykel",
"cykelleasing",
"hyrcykel",
"cykeluthyrning"
],
"amenity/bicycle_repair_station":[
"kedjebrytare",
"Station för cykelreparation",
"cykel",
"tryckluft",
"cykelpump",
"pumpstation",
"cykelreparation"
],
"amenity/biergarten":[
"ölträdgård",
"biergarten",
"servering",
"trädgårdsbar",
"sprit",
"krog",
"utepub",
"utecafé",
"bar",
"Ölträdgård",
"utebar",
"öl",
"pub",
"trädgårdspub",
"uteservering",
"ölcafé"
],
"amenity/binoculars":[
"utsikt",
"Fast monterad kikare",
"kikare",
"fast monterad kikare",
"teleskop"
],
"amenity/boat_rental":[
"båtleasing",
"lånebåt",
"hyrbåt",
"Båtuthyrning",
"båtlån",
"båtuthyrning"
],
"amenity/boat_storage":[
"båt",
"marina",
"båtuppställning",
"uppställning",
"Båtförvaring",
"båthus",
"torrdocka",
"båtförvaring"
],
"amenity/bureau_de_change":[
"växlingskontor",
"resecheckar",
"valuta",
"pengaväxlare",
"pengaväxling",
"Växlingskontor",
"växling",
"pengar"
],
"amenity/bus_station":[
"Busstation / Bussterminal"
],
"amenity/cafe":[
"te",
"kondis",
"kaffeservering",
"servering",
"kaffestuga",
"kafeteria",
"fik",
"cafeteria",
"konditori",
"bistro",
"kaffe",
"Café"
],
"amenity/cafe/bubble_tea":[
"bubbelte",
"taiwanesiskt te",
"boba",
"Bubble tea-café",
"bubble tea-café",
"café. bubble tea"
],
"amenity/cafe/coffee_shop":[
"kaffehus",
"espresso",
"cappuccino",
"americano",
"café",
"varma drycker",
"latte",
"te",
"kakao",
"kaffeaffär",
"Kaffehus",
"bryggkaffe",
"kaffe",
"kaffeshop",
"macchiato"
],
"amenity/car_pooling":[
"bilpoolstation",
"bildelning",
"lånebil",
"hyrbil",
"bilpool",
"Bilpoolstation"
],
"amenity/car_rental":[
"Biluthyrning",
"lånebil",
"hyrbil",
"biluthyrning",
"billån",
"billeasing"
],
"amenity/car_sharing":[
"Bildelningsstation",
"bildelning",
"lånebil",
"hyrbil",
"bilpool",
"bildelningsstation"
],
"amenity/car_wash":[
"biltvätt",
"biltvättanläggning",
"tvättgata",
"tvätt-tunnel",
"portaltvätt",
"Biltvätt"
],
"amenity/casino":[
"spelsalong",
"Kasino",
"poker",
"spelklubb",
"casino",
"spelhåla",
"spelrum",
"tärning",
"blackjack",
"kasino",
"spelhus",
"spel",
"roulette",
"kortspel",
"hasardspel"
],
"amenity/charging_station":[
"snabbladdning",
"laddstation",
"eluttag",
"el",
"Laddstation",
"elbil"
],
"amenity/childcare":[
"dagmamma",
"lekgrupp",
"barnomsorg",
"barnhem",
"dagis",
"Barnomsorg",
"daghem",
"förskola"
],
"amenity/cinema":[
"biograf",
"bioduk",
"biografteater",
"bio",
"film",
"Biograf",
"drive-in"
],
"amenity/clinic":[
"klinik",
"sjukvård",
"distriktssköterska",
"doktor",
"vårdcentral",
"distriktsläkare",
"sjukhus",
"Vårdcentral",
"primärvård",
"läkare"
],
"amenity/clinic/abortion":[
"framkallat missfall",
"abort",
"Abortklinik",
"missfall",
"abortklinik",
"fosterfördrivning",
"avbrytande av havandeskap"
],
"amenity/clinic/fertility":[
"äggfrys",
"barnlöshet",
"fortplantning",
"fertilitetscentrum",
"ägglossning",
"spermie",
"spermadonation",
"fertilitet",
"insemination",
"befruktning",
"reproduktion",
"ivf",
"äggdonation",
"Fertilitetsklinik",
"fertilitetsklinik"
],
"amenity/clock":[
"väggur",
"urtavla",
"kyrkklocka",
"solur",
"klocka",
"Klocka",
"ur",
"väggklocka",
"tidur"
],
"amenity/clock/sundial":[
"gnomon",
"skugga",
"soltid",
"skuggklocka",
"solur",
"solklocka",
"Solur",
"solvisare"
],
"amenity/college":[
"college",
"gymnasium",
"gymnasieområde",
"gymnasie",
"vidareutbildning",
"gymnasiumområde",
"Collegeområde"
],
"amenity/community_centre":[
"folkets hus",
"hembygdsgård",
"bygdegård",
"byalag",
"samlingslokal",
"folkets park",
"byförening",
"Samlingslokal",
"festlokal",
"sockenstuga",
"bystuga",
"evenemang"
],
"amenity/community_centre/lgbtq":[
"hbtq-festlokal",
"hbtq-samlingslokal",
"hbtq--evenemang",
"hbtq",
"HBTQ-samlingslokal"
],
"amenity/compressed_air":[
"Tryckluft",
"tryckluft",
"pumpstation",
"komprimerad luft"
],
"amenity/conference_centre":[
"föreläsning",
"auditorium",
"mässcenter",
"kongresscenter",
"mässa",
"kongresshall",
"utställning",
"Kongresscenter",
"konferens",
"mässhall"
],
"amenity/courthouse":[
"lag",
"rätt",
"juridik",
"Domstol",
"ting",
"rättskipare",
"tribunal",
"instans",
"lagbok",
"domstol"
],
"amenity/coworking_space":[
"Dagkontor"
],
"amenity/crematorium":[
"begravning",
"krematorium",
"Krematorium",
"kremering"
],
"amenity/dentist":[
"tänder",
"tanddoktor",
"tandläkare",
"odontolog",
"tandborstning",
"tand",
"Tandläkare",
"tandhygien",
"tandhygienist"
],
"amenity/dive_centre":[
"sportdykare",
"sportdykning",
"dykare",
"Dykcenter",
"scuba",
"dykning",
"dykcenter",
"grodman"
],
"amenity/doctors":[
"klinik",
"sjukvård",
"sjukvårdare",
"doktor",
"vårdcentral",
"sjukhus",
"läkare",
"vårdinrättning",
"Doktor"
],
"amenity/dojo":[
"kampsport",
"budo",
"japan",
"japansk konst",
"Dojo / Akademi för kampsport",
"kampkonst",
"dojang",
"träningslokal",
"dojo"
],
"amenity/dressing_room":[
"omklädningsrum",
"påklädningsrum",
"loge",
"avklädningsrum",
"påklädning",
"avklädning",
"Omklädningsrum",
"omklädning",
"ombyte"
],
"amenity/drinking_water":[
"dricksvatten",
"källa",
"Dricksvatten",
"fontän",
"vatten"
],
"amenity/driving_school":[
"trafikskola",
"bilskola",
"körkort",
"uppkörning",
"lastbilskort",
"Trafikskola",
"övningskörning",
"körskola"
],
"amenity/embassy":[
"Ambassad"
],
"amenity/events_venue":[
"Evenemangsplats/festlokal",
"dop",
"möten",
"konfirmation",
"festlokal",
"bankettsal",
"fest",
"bröllop",
"festplats",
"möteslokal",
"evenemangsplats",
"konferens",
"födelsedag",
"evenemangslokal"
],
"amenity/exhibition_centre":[
"mässa",
"utställning",
"utställningscenter",
"expo",
"Utställningscenter/Mässa"
],
"amenity/fast_food":[
"skräpmat",
"gatuköksmat",
"hämtmat",
"Snabbmat",
"gatukök",
"snabbmat",
"restaurang",
"takeaway",
"bukfylla",
"junk-food"
],
"amenity/fast_food/burger":[
"mat",
"lunch",
"gatukök",
"restaurang",
"burgare",
"takeaway",
"bukfylla",
"junk-food",
"skräpmat",
"gatuköksmat",
"hämtmat",
"äta",
"snabbmat",
"hamburgare",
"Snabbmat – Hamburgare",
"drive-in",
"grill"
],
"amenity/fast_food/chicken":[
"mat",
"Snabbmat – Kyckling",
"lunch",
"gatukök",
"restaurang",
"takeaway",
"bukfylla",
"junk-food",
"skräpmat",
"gatuköksmat",
"hämtmat",
"äta",
"snabbmat",
"kyckling",
"drive-in",
"grill"
],
"amenity/fast_food/donut":[
"mat",
"gatukök",
"frukost",
"restaurang",
"takeaway",
"bukfylla",
"junk-food",
"café",
"skräpmat",
"gatuköksmat",
"hämtmat",
"äta",
"munkar",
"munk",
"brunch",
"snabbmat",
"donut",
"drive-in",
"kaffe",
"Snabbmat – Munkar"
],
"amenity/fast_food/fish_and_chips":[
"mat",
"lunch",
"fisk och chips",
"gatukök",
"restaurang",
"Snabbmat – Fish & Chips",
"fish and chips",
"takeaway",
"bukfylla",
"junk-food",
"skräpmat",
"gatuköksmat",
"hämtmat",
"äta",
"fish & chips",
"snabbmat",
"drive-in",
"grill"
],
"amenity/fast_food/hot_dog":[
"korvbröd",
"Snabbmat – Korv med bröd",
"snabbmat",
"korv",
"korv med bröd",
"varmkorv"
],
"amenity/fast_food/ice_cream":[
"Snabbmat – Glass"
],
"amenity/fast_food/juice":[
"frukt",
"mat",
"lunch",
"gatukök",
"dryck",
"smoothies",
"fruktdryck",
"shakes",
"Snabbmat – Juice",
"restaurang",
"juice",
"takeaway",
"bukfylla",
"junk-food",
"skräpmat",
"gatuköksmat",
"hämtmat",
"äta",
"snabbmat",
"juicebar",
"drive-in",
"grill"
],
"amenity/fast_food/kebab":[
"mat",
"lunch",
"gatukök",
"restaurang",
"takeaway",
"bukfylla",
"junk-food",
"skräpmat",
"gatuköksmat",
"hämtmat",
"äta",
"snabbmat",
"kebab",
"Snabbmat – Kebab",
"drive-in",
"grill"
],
"amenity/fast_food/mexican":[
"mat",
"lunch",
"gatukök",
"restaurang",
"mexikanskt",
"takeaway",
"bukfylla",
"junk-food",
"skräpmat",
"gatuköksmat",
"hämtmat",
"äta",
"mexico",
"Snabbmat – Mexikanskt",
"snabbmat",
"drive-in",
"grill"
],
"amenity/fast_food/pizza":[
"mat",
"Snabbmat – Pizza",
"lunch",
"pan pizza",
"gatukök",
"restaurang",
"takeaway",
"bukfylla",
"junk-food",
"skräpmat",
"gatuköksmat",
"hämtmat",
"äta",
"pizza",
"pizzeria",
"snabbmat",
"drive-in",
"grill"
],
"amenity/fast_food/sandwich":[
"lunch",
"smörgåsar",
"macka",
"bargetter",
"Snabbmat – Smörgås",
"skräpmat",
"gatuköksmat",
"hämtmat",
"äta",
"smörgås",
"baguetter",
"snabbmat",
"mackor",
"drive-in",
"baguette",
"mat",
"gatukök",
"restaurang",
"takeaway",
"bukfylla",
"junk-food",
"bargett",
"fralla",
"frallor",
"grill"
],
"amenity/ferry_terminal":[
"Färjeterminal"
],
"amenity/fire_station":[
"brandstång",
"brandbil",
"räddningstjänsten",
"brandstation",
"Brandstation",
"brandtorn"
],
"amenity/food_court":[
"mat",
"gatukök",
"mattorg",
"restaurangtorg",
"snabbmat",
"food court",
"restaurang",
"Restaurangtorg"
],
"amenity/fountain":[
"springbrunn",
"fontän",
"Fontän",
"vattenkonst"
],
"amenity/fuel":[
"bensin",
"diesel",
"lng",
"bensinstation",
"Bensinstation",
"bränsle",
"propan",
"tapp",
"tankstation",
"cng",
"mack",
"biodiesel"
],
"amenity/gambling":[
"spelhall",
"poker",
"casino",
"keno",
"vadslagning",
"Spelhall",
"blackjack",
"kasino",
"spel",
"slots",
"roulette",
"spelautomater",
"bingo",
"lotteri"
],
"amenity/give_box":[
"donering",
"free box",
"skänka bort",
"frilåda",
"donation",
"free table",
"bortskänkningslåda",
"fritt bord",
"Bortskänkningslåda"
],
"amenity/grave_yard":[
"urnlund",
"gravplats",
"griftegård",
"kyrkogård",
"begravningsplats",
"Kyrkogård",
"minneslund"
],
"amenity/grit_bin":[
"sand",
"salt",
"sandlåda",
"halkbekämpning",
"Sandkista",
"sandkista",
"sandbehållare",
"halka"
],
"amenity/hospital":[
"sanatorium",
"sjukhus",
"läkare",
"sjukhusområde",
"Sjukhusområde",
"klinik",
"sjukvård",
"institution",
"lasarett",
"läkarmottagning",
"sjukstuga",
"vårdhem",
"kirurgi",
"sjuk"
],
"amenity/hunting_stand":[
"jakt",
"skjuta",
"viltjakt",
"Jakttorn",
"utkik",
"skjutstege",
"älgtorn",
"utkikstorn",
"vilt",
"jakttorn"
],
"amenity/ice_cream":[
"glasskiosk",
"yogurt",
"glass",
"Glassaffär",
"mjukglass",
"sorbet",
"sherbet",
"frozen",
"kulglass",
"gelato",
"glassaffär"
],
"amenity/internet_cafe":[
"internetkafé",
"internetcafé",
"internetcaffe",
"internetcafe",
"cybercafé",
"Internetkafé"
],
"amenity/karaoke_box":[
"karaoke box",
"karaoke-rum",
"karaoke-tv",
"karaoke-klubb",
"Karaoke Box",
"ktv",
"karaoke lounge"
],
"amenity/kindergarten":[
"kindergarten",
"lekplats",
"Förskoleområde",
"dagis",
"lekskola",
"daghem",
"lekis",
"förskola"
],
"amenity/kneipp_water_cure":[
"kallvattenkuranstalt",
"vattenkur",
"kallvattenkur",
"kneipp vattenterapi",
"kneipp",
"hydrotherapie",
"Kneipp vattenterapi",
"fotbad. vatten"
],
"amenity/language_school":[
"språk",
"språkskola",
"språkkurs",
"Språkskola",
"språkutbildning",
"esl"
],
"amenity/lavoir":[
"tvättstuga",
"tvättning",
"tvättställe",
"Tvättbrygga",
"klädtvätt",
"tvättbrygga",
"tvätt",
"lavoir",
"kläder",
"handtvätt"
],
"amenity/letter_box":[
"Postlåda",
"brevlåda",
"brevinkast",
"postlucka",
"postlåda"
],
"amenity/library":[
"läsesal",
"bibliotek",
"bokrum",
"Bibliotek",
"boksamling",
"bibbla",
"böcker",
"bokskatt",
"bok"
],
"amenity/loading_dock":[
"lager",
"lastbrygga",
"dörr",
"lastning",
"lagerhus",
"Lastkaj",
"gods",
"utlastning",
"inlastning",
"fraktbrygga",
"frakt",
"lastkaj"
],
"amenity/lounger":[
"soldäck",
"solning",
"Solstol(ar)",
"solstolar",
"stolar",
"bänkar"
],
"amenity/love_hotel":[
"kärlekshotell",
"Kärlekshotell",
"hotell",
"sexhotell",
"korttidshotell"
],
"amenity/marketplace":[
"saluhall",
"Marknadsplats",
"salutorg",
"marknad",
"torg"
],
"amenity/monastery":[
"helgedom",
"allah",
"församling",
"tempelområde",
"kyrka",
"katedral",
"religiös anläggning",
"kor",
"vallfärdsort",
"andaktsrum",
"gudshus",
"tillbedjan",
"moské",
"begravningskapell",
"andligt område",
"moske",
"fristad",
"kloster",
"dopkapell",
"kapell",
"gudstjänstslokal",
"tro",
"mission",
"bönehus",
"gud",
"dyrkan",
"guds hus",
"kristendom",
"missionshus",
"sanktuarium",
"andaktssal",
"dom",
"kyrkogård",
"böneplats",
"basilika",
"tempel",
"kyrkobyggnad",
"religiös",
"religiöst område",
"Klosterområde",
"bönhus",
"sidokapell",
"kranskapell",
"predikan",
"vallfärgsplats",
"betel",
"kristen",
"kyrkbyggnad",
"synagoga",
"mässkapell",
"religion",
"annexkyrka",
"gravkapell",
"kyrkorum",
"andaktslokal",
"gudstjänstlokal",
"gudstjänst",
"kyrksal",
"korkapell",
"tabernakel"
],
"amenity/money_transfer":[
"finans",
"räkning",
"valuta",
"utbetalning",
"pengaöverföring",
"betalning",
"inbetalning",
"Pengaöverföring",
"valutaöverföring",
"faktura",
"kontanter",
"pengar"
],
"amenity/mortuary":[
"minneshem",
"död",
"krematorium",
"Bårhus",
"likförvaring",
"bårhus",
"likbod",
"begravningsplats",
"begravningsbyrå",
"lik"
],
"amenity/motorcycle_parking":[
"motorcykelställ",
"parkeringsplats",
"motorcykelparkering",
"ställplats",
"motorcykel",
"parkering motorcykel",
"parkeringsplats motorcykel",
"parkering",
"Motorcykelparkering"
],
"amenity/motorcycle_rental":[
"motorcykeluthyrning",
"minibike",
"hyrmotorcykel",
"motorcykelleasing",
"motorcykel",
"moped",
"dirt bike",
"scooter",
"Motorcykeluthyrning",
"sidovagn",
"motorscooter",
"motorcykellån"
],
"amenity/music_school":[
"musikskola",
"musikinstrument",
"sångskola",
"kultur",
"kör",
"instrument",
"musik",
"kulturskola",
"instrumentskola",
"sång",
"Musikskola"
],
"amenity/nightclub":[
"diskotek",
"dansställe",
"klubb",
"bar",
"nattklubb",
"nöjeslokal",
"Nattklubb",
"disco",
"disko*",
"dans",
"dansklubb"
],
"amenity/nightclub/lgbtq":[
"lesbisk klubb",
"HBTQ-nattklubb",
"gay nattklub",
"hbtq-nattklubb",
"lesbisk nattklubb",
"lesbiskt disko",
"gay disko",
"gay-klubb",
"gay-nattklubb",
"gay-disko",
"hbtq-klubb"
],
"amenity/nursing_home":[
"Vårdhem"
],
"amenity/parking":[
"parkeringsplats",
"bil",
"p-plats",
"bilparkering",
"parkeringsområde",
"Parkeringsplats",
"parkering"
],
"amenity/parking/multi-storey":[
"parkeringsbyggnad",
"flervånig",
"bil",
"flervånig parkeringsgarage",
"parkeringshus",
"garage",
"bilparkering",
"parkeringsgarage",
"inomhusparkering",
"flervånig bilparkering",
"parkering",
"parkeringsramp",
"parkeringsdäck",
"garagebyggnad",
"Flervånigt parkeringsgarage"
],
"amenity/parking/park_ride":[
"pendling",
"parkeringsplats",
"bil",
"infartsparkering",
"p-plats",
"bilparkering",
"parkeringsområde",
"pendelparkeringsplats",
"parkering",
"Pendelparkeringsplats",
"pendlare",
"pendelparkering",
"pendlarparkering"
],
"amenity/parking/underground":[
"underjordisk parkering",
"parkeringsplats",
"fordonsparkering",
"Underjordisk parkering",
"p-plats",
"bilparkering",
"parkeringshus",
"parkeringsgarage",
"parkeringsområde",
"underjordisk",
"parkering"
],
"amenity/parking_entrance":[
"utfart",
"garage",
"parkeringshus",
"infart",
"parkeringsgarage",
"In- och utfart parkeringsgarage"
],
"amenity/parking_space":[
"parkeringsruta",
"handikapsparkering",
"handikapsficka",
"Parkeringsruta",
"enskild parkeringsplats",
"parkeringsyta",
"parkeringsficka"
],
"amenity/parking_space/disabled":[
"handikapad",
"handikappsplats",
"rullstolsplats",
"rullstol",
"handikapsparkering",
"Handikappsplats",
"handikapsficka"
],
"amenity/payment_centre":[
"räkning",
"valuta",
"utbetalning",
"betalningskontor",
"inbetalning",
"check",
"kontanter",
"skatt",
"betalning",
"betalningscenter",
"faktura",
"pengar",
"Betalningscenter"
],
"amenity/payment_terminal":[
"Betalningsterminal",
"räkning",
"valuta",
"överföring",
"betalningsterminal",
"utbetalning",
"inbetalning",
"ekiosk",
"kontanter",
"skatteinbetalning",
"skatt",
"betalning",
"pengaröverföring",
"atm",
"faktura",
"pengar"
],
"amenity/pharmacy":[
"Läkemedel",
"drog*",
"medicin",
"läkemedel*",
"droghandel",
"apotek",
"läkemedelsaffär",
"farmaceut",
"recept"
],
"amenity/photo_booth":[
"fotobås",
"bild",
"Fotoautomat",
"foto",
"kameraautomat",
"fotoautomat",
"kamera"
],
"amenity/place_of_worship":[
"helgedom",
"allah",
"församling",
"tempelområde",
"kyrka",
"katedral",
"religiös anläggning",
"kor",
"vallfärdsort",
"andaktsrum",
"gudshus",
"tillbedjan",
"moské",
"begravningskapell",
"andligt område",
"moske",
"fristad",
"kloster",
"dopkapell",
"kapell",
"gudstjänstslokal",
"tro",
"mission",
"bönehus",
"gud",
"dyrkan",
"guds hus",
"kristendom",
"missionshus",
"sanktuarium",
"andaktssal",
"dom",
"kyrkogård",
"böneplats",
"basilika",
"tempel",
"kyrkobyggnad",
"religiös",
"religiöst område",
"Plats för tillbedjan",
"bönhus",
"sidokapell",
"kranskapell",
"socken",
"predikan",
"vallfärgsplats",
"betel",
"kristen",
"kyrkbyggnad",
"synagoga",
"mässkapell",
"religion",
"slottskapell",
"annexkyrka",
"gravkapell",
"kyrkorum",
"andaktslokal",
"gudstjänstlokal",
"gudstjänst",
"kyrksal",
"korkapell",
"pastorat",
"tabernakel"
],
"amenity/place_of_worship/buddhist":[
"pagoda",
"Buddhisttempel",
"kloster",
"buddha",
"meditation",
"zendo",
"buddhism",
"chörten",
"stupa",
"tempel",
"dojo",
"vihara"
],
"amenity/place_of_worship/christian":[
"helgedom",
"församling",
"tempelområde",
"kyrka",
"katedral",
"religiös anläggning",
"kor",
"vallfärdsort",
"andaktsrum",
"gudshus",
"tillbedjan",
"begravningskapell",
"andligt område",
"fristad",
"kloster",
"dopkapell",
"kapell",
"gudstjänstslokal",
"tro",
"mission",
"bönehus",
"gud",
"dyrkan",
"guds hus",
"kristendom",
"missionshus",
"sanktuarium",
"Kristen kyrka",
"andaktssal",
"dom",
"kyrkogård",
"böneplats",
"basilika",
"tempel",
"kyrkobyggnad",
"religiös",
"religiöst område",
"bönhus",
"sidokapell",
"kranskapell",
"socken",
"predikan",
"vallfärgsplats",
"betel",
"kristen",
"kyrkbyggnad",
"mässkapell",
"religion",
"slottskapell",
"annexkyrka",
"gravkapell",
"kyrkorum",
"andaktslokal",
"gudstjänstlokal",
"gudstjänst",
"kyrksal",
"korkapell",
"pastorat",
"tabernakel"
],
"amenity/place_of_worship/christian/jehovahs_witness":[
"bönehus",
"Rikets sal för Jehovas vittne",
"kyrka",
"hus för tillbedjan",
"jehovas vittne",
"guds hus",
"rikets sal för jehovas vittne",
"tillbedjan",
"bön",
"kristen",
"rikets sal",
"kristendom"
],
"amenity/place_of_worship/christian/la_luz_del_mundo":[
"bönehus",
"världens ljuskyrka",
"hus för bön",
"kyrka",
"guds hus",
"la luz del mundo-tempel",
"kristen",
"the light of the world-kyrka",
"La Luz del Mundo-tempel",
"kristendom",
"la luz del mundo",
"tempel"
],
"amenity/place_of_worship/christian/quaker":[
"kväkarevännernas möteshus",
"bönehus",
"hus för bön",
"kväkare",
"guds hus",
"Kväkarevännernas möteshus",
"kristen",
"kristendom",
"vännernas samfund"
],
"amenity/place_of_worship/hindu":[
"hinduism",
"sanatana dharma",
"helgedom",
"hindu",
"Hindutempel",
"garbhagriha",
"puja",
"arcana",
"tempel"
],
"amenity/place_of_worship/jewish":[
"helgedom",
"dom",
"predikan",
"judisk",
"katedral",
"synagoga",
"böneplats",
"tempel",
"religion",
"tro",
"bönehus",
"Judisk synagoga",
"gudshus",
"gudstjänstlokal",
"tillbedjan",
"jude",
"judendom",
"missionshus"
],
"amenity/place_of_worship/muslim":[
"helgedom",
"muslim",
"muslimsk",
"predikan",
"böneplats",
"religion",
"kyrkobyggnad",
"tro",
"bönehus",
"gudshus",
"gudstjänstlokal",
"Muslimsk moské",
"tillbedjan",
"moské",
"minaret"
],
"amenity/place_of_worship/shinto":[
"kami",
"helgedom",
"jinja",
"torii",
"shintohelgedom",
"shrine",
"tempel",
"yashiro",
"jingū",
"shinto shrine",
"miya",
"Jinja (Shintoistisk helgedom)",
"shintoism",
"shinto"
],
"amenity/place_of_worship/sikh":[
"helgedom",
"gurudwara",
"sikh",
"Sikhiskt tempel",
"sikhtempel",
"sikh-tempel",
"sikhism",
"tempel"
],
"amenity/place_of_worship/taoist":[
"helgedom",
"Taoistiskt tempel",
"tao",
"taoism",
"taoistiskt tempel",
"daoism",
"tempel"
],
"amenity/planetarium":[
"museum",
"planetarium",
"observatorium",
"astronomi",
"Planetarium"
],
"amenity/police":[
"polisman",
"pass",
"poliskonstapel",
"polis",
"Polis",
"snut",
"polismyndighet",
"kriminalare",
"ordningsmakt",
"polisväsende",
"lag",
"konstapel",
"polismakt",
"polisstation"
],
"amenity/polling_station":[
"val",
"rösta",
"omröstning",
"röstmaskin",
"vallokal",
"valbås",
"valsedel",
"röstning",
"folkomröstning",
"valmaskin",
"valurna",
"omröstningsapparat",
"Permanent vallokal"
],
"amenity/post_box":[
"brevlåda",
"brevinlämning",
"brevinkast",
"postfack",
"post",
"postbox",
"Brevlåda",
"paketinlämning",
"postlåda",
"brev"
],
"amenity/post_depot":[
"brevsortering",
"post",
"postsorteringskontor",
"postterminal",
"postdistribution",
"sortering",
"Postsorteringskontor",
"postsortering",
"brev",
"brevdistribution"
],
"amenity/post_office":[
"Postkontor",
"postkontor",
"post",
"kort",
"postverk",
"posten",
"frimärke",
"paket",
"försändelser",
"postgång",
"postväsende",
"brev"
],
"amenity/prep_school":[
"kvälsskola",
"matematik",
"akademisk",
"testförberedelse",
"Pluggskola",
"läxa",
"läsning",
"pluggskola",
"läxhjälp",
"handledning",
"skrivning"
],
"amenity/prison":[
"häkte",
"fångvårdsanstalt",
"polisarrest",
"fängelse",
"arrest",
"Fängelseområde",
"anstalt",
"fängelseförvar",
"fängelseområde",
"fånganstalt",
"finka"
],
"amenity/pub":[
"bar",
"ölservering",
"nattklubb",
"öl",
"sprit",
"alkohol",
"ölstuga",
"drinkar",
"pub",
"Pub",
"krog"
],
"amenity/pub/irish":[
"irland",
"irländsk",
"bar",
"irländsk bar",
"irländsk pub",
"pub",
"Irländsk pub"
],
"amenity/pub/lgbtq":[
"lesbisk pub",
"lgbtq pub",
"lgbt pub",
"HBTQ-pub",
"gay-pub",
"hbtq-pub",
"lgb pub"
],
"amenity/pub/microbrewery":[
"ölframställning",
"brewpub",
"alkohol",
"sprit",
"öltillverkning",
"drink",
"Brewpub",
"mikrobryggeri",
"bar",
"öl",
"bryggeri",
"pub",
"hantverksbryggeri"
],
"amenity/public_bath":[
"badinrättning",
"het källa",
"badhus",
"simbassäng",
"bad",
"bassängbad",
"bassäng",
"badplats",
"publikt bad",
"strandbad",
"onsen",
"strand",
"Publikt bad",
"fotbad",
"badställe"
],
"amenity/public_bookcase":[
"begagnade böcker",
"publik bokhylla",
"Offentlig bokhylla",
"låneböcker",
"bokdelning",
"bibliotek",
"offentlig bokhylla",
"bokbyte"
],
"amenity/ranger_station":[
"informationscenter",
"infocenter",
"besökscenter",
"friluftsanläggningen",
"friluftsområde",
"park",
"friluftsliv",
"Friluftsanläggningen"
],
"amenity/recycling":[
"Återvinning"
],
"amenity/recycling/container/electrical_items":[
"elektronikskrot",
"surfplattor",
"återvinningsstation",
"Elektronikskrot",
"elektronik",
"datorer",
"elektroniskt avfall",
"elektronikåtervinning",
"telefoner",
"återbruk",
"återvinning",
"elskrot"
],
"amenity/recycling/container/green_waste":[
"kompost",
"skräp",
"biologiskt nedbrytbart",
"biologiskt",
"komposterbart",
"nedbrytbart",
"Komposterbart",
"trädgårdsavfall",
"matavfall",
"organiskt",
"trädgård",
"sopor"
],
"amenity/recycling_centre":[
"skräp",
"återvinningsstation",
"flaskor",
"dumpa",
"Återvinningscentral",
"glas",
"sopstation",
"skrot",
"återbruk",
"burkar",
"återvinning",
"sopor"
],
"amenity/recycling_container":[
"skräp",
"container",
"metall",
"Återvinningscontainer",
"återvinningscontainer",
"återvinningsstation",
"flaskor",
"glas",
"återbruk",
"sopstation",
"skrot",
"burkar",
"återvinning",
"sopor"
],
"amenity/refugee_site":[
"flykting",
"flyktingläger",
"evakueringsläger",
"migranter",
"flyktingar",
"Flyktingläger"
],
"amenity/research_institute":[
"forskningslaboratorium",
"forskningsinstitutsområde",
"experiment",
"forskning",
"tillämpad forskning",
"forskningsinstitution",
"forskningslaboratorier",
"institut",
"forskning och utveckling",
"Forskningsinstitutsområde",
"forskningsinstitut",
"fou"
],
"amenity/restaurant":[
"café. matsal",
"lunch",
"servering",
"grillbar",
"värdshus",
"restaurang",
"kafé",
"brasserie",
"cafeteria",
"krog",
"bodega",
"rotisseri",
"matservering",
"bar",
"matställe",
"pizzeria",
"restauration",
"pub",
"Restaurang",
"näringsställe",
"sylta",
"kaffe"
],
"amenity/restaurant/american":[
"lunch",
"usa",
"servering",
"grillbar",
"värdshus",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"matställe",
"näringsställe",
"kaffe",
"café. matsal",
"restaurang",
"kafé",
"amerikansk mat",
"bodega",
"rotisseri",
"pizzeria",
"restauration",
"pub",
"amerikansk restaurang",
"sylta",
"Amerikansk restaurang"
],
"amenity/restaurant/asian":[
"café. matsal",
"asiatisk restaurang",
"lunch",
"servering",
"grillbar",
"värdshus",
"restaurang",
"kafé",
"brasserie",
"cafeteria",
"krog",
"bodega",
"rotisseri",
"matservering",
"bar",
"matställe",
"Asiatisk restaurang",
"pizzeria",
"asiatisk mat",
"restauration",
"pub",
"näringsställe",
"sylta",
"kaffe"
],
"amenity/restaurant/chinese":[
"lunch",
"servering",
"grillbar",
"värdshus",
"kinesisk",
"kinesisk restaurang",
"brasserie",
"cafeteria",
"kinamat",
"krog",
"matservering",
"bar",
"Kinesisk restaurang",
"matställe",
"näringsställe",
"kaffe",
"café. matsal",
"kina",
"restaurang",
"kafé",
"bodega",
"rotisseri",
"pizzeria",
"restauration",
"pub",
"sylta"
],
"amenity/restaurant/french":[
"fransk restaurang",
"lunch",
"servering",
"grillbar",
"värdshus",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"matställe",
"Fransk restaurang",
"näringsställe",
"kaffe",
"café. matsal",
"restaurang",
"kafé",
"bodega",
"rotisseri",
"pizzeria",
"frankrike",
"restauration",
"pub",
"fransk mat",
"sylta"
],
"amenity/restaurant/german":[
"lunch",
"servering",
"grillbar",
"värdshus",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"matställe",
"tysk mat",
"näringsställe",
"kaffe",
"tysk restaurang",
"café. matsal",
"tyskland",
"restaurang",
"kafé",
"Tysk restaurang",
"bodega",
"rotisseri",
"pizzeria",
"restauration",
"pub",
"sylta"
],
"amenity/restaurant/greek":[
"Grekisk restaurang",
"lunch",
"servering",
"grillbar",
"värdshus",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"matställe",
"grekisk restaurang",
"näringsställe",
"kaffe",
"café. matsal",
"grekisk mat",
"restaurang",
"kafé",
"bodega",
"rotisseri",
"grekland",
"pizzeria",
"restauration",
"pub",
"sylta"
],
"amenity/restaurant/indian":[
"lunch",
"servering",
"grillbar",
"värdshus",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"matställe",
"indisk restaurang",
"näringsställe",
"kaffe",
"indisk mat",
"café. matsal",
"restaurang",
"kafé",
"bodega",
"rotisseri",
"pizzeria",
"Indisk restaurang",
"indien",
"restauration",
"pub",
"sylta"
],
"amenity/restaurant/italian":[
"lunch",
"servering",
"grillbar",
"värdshus",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"matställe",
"Italiensk restaurang",
"italien",
"näringsställe",
"kaffe",
"café. matsal",
"restaurang",
"kafé",
"bodega",
"rotisseri",
"italiensk mat",
"pizzeria",
"restauration",
"pub",
"sylta",
"italiensk restaurang"
],
"amenity/restaurant/japanese":[
"lunch",
"servering",
"Japansk restaurang",
"grillbar",
"värdshus",
"japan",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"matställe",
"näringsställe",
"kaffe",
"café. matsal",
"japansk restaurang",
"restaurang",
"kafé",
"bodega",
"rotisseri",
"pizzeria",
"japansk mat",
"restauration",
"pub",
"sylta"
],
"amenity/restaurant/mexican":[
"lunch",
"servering",
"grillbar",
"värdshus",
"mexikansk restaurang",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"matställe",
"näringsställe",
"kaffe",
"café. matsal",
"Mexikansk restaurang",
"restaurang",
"mexiko",
"kafé",
"bodega",
"rotisseri",
"pizzeria",
"mexikansk mat",
"restauration",
"pub",
"sylta"
],
"amenity/restaurant/noodle":[
"lunch",
"servering",
"grillbar",
"värdshus",
"risnudlar",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"matställe",
"nudlar",
"ris",
"näringsställe",
"kaffe",
"café. matsal",
"Nudelrestaurang",
"restaurang",
"kafé",
"nudelrestaurang",
"bodega",
"rotisseri",
"pizzeria",
"restauration",
"pub",
"sylta"
],
"amenity/restaurant/pizza":[
"lunch",
"servering",
"grillbar",
"värdshus",
"brasserie",
"cafeteria",
"krog",
"pan-pizza",
"matservering",
"bar",
"matställe",
"pizza",
"panpizza",
"näringsställe",
"kaffe",
"café. matsal",
"pan pizza",
"restaurang",
"pizzarestaurang",
"kafé",
"bodega",
"rotisseri",
"pizzeria",
"restauration",
"pub",
"Pizzarestaurang",
"sylta"
],
"amenity/restaurant/seafood":[
"hummer",
"lunch",
"kräftdjur",
"servering",
"grillbar",
"värdshus",
"blötdjur",
"Fisk- och skaldjursrestaurang",
"brasserie",
"cafeteria",
"krog",
"krabba",
"fiskerestaurang",
"matservering",
"bar",
"matställe",
"bläckfisk",
"näringsställe",
"kaffe",
"café. matsal",
"seafood",
"fisk- och skaldjursrestaurang",
"restaurang",
"kafé",
"bodega",
"skaldjur",
"rotisseri",
"räkor",
"skaldjursrestaurang",
"fisk",
"ostron",
"krabbor",
"pizzeria",
"restauration",
"pub",
"sylta",
"musslor"
],
"amenity/restaurant/steakhouse":[
"lunch",
"servering",
"grillbar",
"värdshus",
"steakhouse",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"matställe",
"steak house",
"näringsställe",
"kaffe",
"kött",
"café. matsal",
"Stekhus",
"biff",
"restaurang",
"kafé",
"bodega",
"rotisseri",
"pizzeria",
"restauration",
"pub",
"slakthus",
"sylta",
"stekhus"
],
"amenity/restaurant/sushi":[
"lunch",
"servering",
"grillbar",
"värdshus",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"matställe",
"asiatisk mat",
"sushi",
"näringsställe",
"kaffe",
"sushi-restaurang",
"café. matsal",
"asiatisk restaurang",
"restaurang",
"kafé",
"bodega",
"rotisseri",
"Sushi-restaurang",
"pizzeria",
"restauration",
"pub",
"sylta"
],
"amenity/restaurant/thai":[
"lunch",
"servering",
"grillbar",
"värdshus",
"Thai-restaurang",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"matställe",
"asiatisk mat",
"thai-restaurang",
"thaimat",
"thailand",
"näringsställe",
"kaffe",
"café. matsal",
"asiatisk restaurang",
"restaurang",
"thai",
"kafé",
"bodega",
"rotisseri",
"pizzeria",
"restauration",
"pub",
"sylta"
],
"amenity/restaurant/turkish":[
"lunch",
"turkisk restaurang",
"servering",
"grillbar",
"värdshus",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"matställe",
"näringsställe",
"kaffe",
"café. matsal",
"Turkisk restaurang",
"restaurang",
"kafé",
"turkiet",
"bodega",
"rotisseri",
"turkisk mat",
"turkisk",
"pizzeria",
"restauration",
"pub",
"sylta"
],
"amenity/restaurant/vietnamese":[
"lunch",
"vietnamesisk restaurang",
"servering",
"grillbar",
"värdshus",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"matställe",
"asiatisk mat",
"Vietnamesisk restaurang",
"näringsställe",
"kaffe",
"café. matsal",
"asiatisk restaurang",
"vietnam",
"restaurang",
"kafé",
"bodega",
"rotisseri",
"pizzeria",
"vietnamesisk mat",
"restauration",
"pub",
"sylta"
],
"amenity/sanitary_dump_station":[
"tömningsplats",
"gråvatten",
"toalettömning",
"Latrintömning för campingfordon",
"sanitet",
"latrintömning",
"campingplats",
"torrtoalett",
"campingtoalett"
],
"amenity/school":[
"högskoleområde",
"gymnasium",
"grundskola",
"campus",
"Skolområde",
"skolgård",
"universitet",
"högskola",
"högstadium",
"mellanstadium",
"universitetsområde",
"skolområde",
"lågstadium"
],
"amenity/shelter":[
"väntkur",
"grotta",
"hydda",
"skydd",
"vindskydd",
"Väderskydd",
"koja",
"väderskydd",
"tak över huvudet",
"picknick",
"lusthus"
],
"amenity/shelter/gazebo":[
"trädgårdspaviljong",
"fåfänga",
"paviljong",
"Lusthus",
"kolonistuga",
"lusthus"
],
"amenity/shelter/lean_to":[
"vindskydd",
"gapskjul",
"Vindskydd",
"skärmskydd"
],
"amenity/shelter/picnic_shelter":[
"Picknicktak",
"picknickplats",
"rastplats",
"paviljong",
"pavilion",
"utflykt",
"picknicktak",
"picknick"
],
"amenity/shelter/public_transport":[
"busskur",
"busshållplats",
"väntplats",
"skydd",
"väderskydd för kollektivtrafik",
"väderskydd",
"spårvagnshållplats",
"Väderskydd för kollektivtrafik"
],
"amenity/shower":[
"duschbad",
"Dusch",
"duschrum",
"badrum",
"duschkabin",
"duschutrymme",
"dusch"
],
"amenity/smoking_area":[
"rökruta",
"cigarett",
"Rökområde",
"rökning tillåten",
"rökrum",
"röka",
"rökning",
"rökområde"
],
"amenity/social_centre":[
"musikskola",
"Medborgarhus",
"kurser",
"utbildning",
"kulturskola",
"folkets park",
"möte",
"evenemang",
"fest",
"möteslokal",
"förbund",
"föreningslokal",
"kultur",
"lokal",
"kulturverksamhet",
"nöje",
"förening",
"kurs",
"föreningsgård",
"allaktivitetshus",
"event",
"medborgarhus"
],
"amenity/social_facility":[
"social inrättning",
"uteliggare",
"social",
"välgörenhetsorganisationer",
"social hjälp",
"socialen",
"välgörenhet",
"hjälparbete",
"Social inrättning"
],
"amenity/social_facility/ambulatory_care":[
"öppenvård",
"Öppenvård",
"ambulerande vård",
"vård",
"hemvård",
"hemtjänst"
],
"amenity/social_facility/food_bank":[
"matbank",
"Matbank",
"välgörenhetsorganisation",
"matutdelning",
"matpaket"
],
"amenity/social_facility/group_home":[
"gruppboende",
"grupphem",
"välgörenhetsorganisationer",
"gammal",
"välgörenhet",
"hjälparbete",
"ålderdomshem",
"kollektiv",
"Gruppboende"
],
"amenity/social_facility/homeless_shelter":[
"Härbärge",
"hemlös",
"sovsal",
"härbärge",
"bostadslös"
],
"amenity/social_facility/nursing_home":[
"pensionärshem",
"servicehus",
"hem för gamla",
"Seniorboende",
"servicehem",
"hvb-hem",
"äldreboende",
"seniorboende",
"senior",
"pensionär",
"vårdhem",
"assistansboende",
"ålderdomshem",
"hem för vård och boende"
],
"amenity/studio":[
"studio",
"utsändningslokal",
"tv",
"filminspelning",
"inspelningslokal",
"television",
"inspelning",
"filmstudio",
"radiostudio",
"tv-studio",
"Studio",
"radio"
],
"amenity/studio/audio":[
"inspelningsstudio",
"ljudstudio",
"ljudinspelning",
"ljudproduktion",
"ljudmix",
"Inspelningsstudio",
"sångstudio"
],
"amenity/studio/radio":[
"studio",
"radiosändning",
"sändning",
"fm",
"Radiostation",
"radiostation",
"am",
"radiostudio",
"radio"
],
"amenity/studio/television":[
"studio",
"tv",
"television",
"tv-sändning",
"TV-studio",
"tv-station",
"tv-studio"
],
"amenity/studio/video":[
"filminspelning",
"videoinspelning",
"Filmstudio",
"videoproduktion",
"filmstudio",
"film",
"video",
"filmproduktion"
],
"amenity/taxi":[
"taxificka",
"taxistation",
"taxi",
"taxihållplats",
"Taxihållplats"
],
"amenity/telephone":[
"telefonautomat",
"telefonkiosk",
"telefonkur",
"telefon",
"telefonhytt",
"Telefon"
],
"amenity/theatre":[
"skådebana",
"drama",
"Teater",
"teaterföreställning",
"föreställning",
"skådespel",
"skådeplats",
"scen",
"musikal",
"pjäs",
"teater"
],
"amenity/theatre/type/amphi":[
"utomhus",
"utomhusteater",
"läktare",
"amfiteater",
"scen",
"teater",
"Amfiteater",
"utescen"
],
"amenity/toilets":[
"avträde",
"latrin",
"hemlighus",
"skithus",
"badrum",
"toa",
"Toaletter",
"utedass",
"bekvämlighetsinrättning",
"wc",
"baja-maja",
"klo",
"vattentoalett",
"dass",
"torrklosett",
"klosett",
"toalett",
"vattenklosett",
"bajamaja",
"mugg"
],
"amenity/toilets/disposal/flush":[
"badrum",
"Vattentoalett",
"toalett",
"spoltoalett",
"wc",
"vattentoalett"
],
"amenity/toilets/disposal/pitlatrine":[
"grop-latrin",
"uthus",
"dass",
"toalett",
"Grop-latrin",
"groptoalett"
],
"amenity/toilets/portable":[
"Portabel toalett",
"kemisk toalett",
"mobil toalett",
"toalett",
"bajamaja",
"porta",
"portabel toalett"
],
"amenity/townhall":[
"stadshus",
"ämbetsverk",
"folkets hus",
"fullmäktige",
"riksdag",
"domstolsbyggnad",
"parlament",
"samlingslokal",
"myndighet",
"representation",
"samlingsplats",
"stad",
"Kommunhus",
"kommunalhus",
"by",
"kommun",
"kommunstyrelse",
"förvaltning"
],
"amenity/townhall/city":[
"stadshus",
"kommunhus",
"regering",
"Rådhus",
"borgmästare",
"rådhus",
"kommun",
"tingshus"
],
"amenity/toy_library":[
"spel",
"Leksaksbibliotek",
"leksak",
"leksaksbibliotek"
],
"amenity/university":[
"college",
"universitetsbyggnad",
"högskola",
"högskoleområde",
"universitetsområde",
"akademi",
"universitet",
"Universitetsområde",
"lärosäte"
],
"amenity/vacuum_cleaner":[
"Dammsugarstation",
"bildammsugare",
"sugstation",
"bilsugare",
"bildtvätt",
"dammsugarstation"
],
"amenity/vehicle_inspection":[
"bilprovning",
"Fordonsbesiktning",
"bilprovningen",
"fordonsinspektion",
"besiktning",
"fordonsbesiktning",
"bilbesiktning",
"bilinspektion"
],
"amenity/vending_machine":[
"biljett",
"tuggummiautomater",
"läsk",
"biljettautomat",
"Varuautomat",
"varuautomat",
"läskautomat",
"varumaskin",
"biljetter",
"godisautomat",
"mellanmål"
],
"amenity/vending_machine/bottle_return":[
"pantautomat",
"pantmaskin",
"Pantautomat"
],
"amenity/vending_machine/bread":[
"brödautomat",
"bröd",
"mat",
"matvarumaskin",
"matautomat",
"varuautomat",
"Brödvarumaskin",
"varumaskin",
"matvaruautomat"
],
"amenity/vending_machine/cigarettes":[
"cigarettautomat",
"cigaretter",
"snusautomat",
"tobaksautomat",
"Cigarettautomat"
],
"amenity/vending_machine/coffee":[
"the",
"te",
"kaffeautomat",
"espresso",
"expresso",
"varuautomat",
"Kaffeautomat",
"varumaskin",
"kaffe"
],
"amenity/vending_machine/condoms":[
"kondomomat",
"kondomautomat",
"Kondomautomat",
"kondomer"
],
"amenity/vending_machine/drinks":[
"kaffeautomat",
"drickautomat",
"läsk",
"dryck",
"dryckesautomat",
"läskautomat",
"kaffemaskin",
"juice",
"kaffe",
"Dryckesautomat",
"dryckautomat"
],
"amenity/vending_machine/eggs":[
"äggvarumaskin",
"mat",
"matvarumaskin",
"Äggvarumaskin",
"matautomat",
"ägg",
"varuautomat",
"äggautomat",
"varumaskin",
"matvaruautomat",
"äggmaskin"
],
"amenity/vending_machine/electronics":[
"kabel",
"laddare",
"kablar",
"varumaskin",
"laddkabel",
"laddkablar",
"varumaskin för elektronik",
"mobiltelefon",
"pekplatta",
"telefon",
"surfplatta",
"varuautomat",
"elektronik",
"Varumaskin för elektronik",
"öronsnäckor",
"hörlurar"
],
"amenity/vending_machine/elongated_coin":[
"mynt",
"minnesmyntmaskin",
"elongated penny",
"myntpressmaskin",
"ecm",
"coin maskin",
"minne",
"minnesmynt",
"penny press",
"souvenirmynt",
"elongated coin-maskin",
"Elongated coin-maskin (myntpressmaskin)",
"elongated coin",
"souvenir"
],
"amenity/vending_machine/excrement_bags":[
"hundpåsar",
"hund",
"bajs",
"hundskit",
"Bajspåsar",
"hundbajs",
"avföringspåse",
"djur",
"bajspåsar",
"skitpåse",
"hundbajspåsar"
],
"amenity/vending_machine/feminine_hygiene":[
"kvinnor",
"Varumaskin för mensskydd",
"varumaskin för mensskydd",
"binda",
"tampong",
"kvinna",
"bindor",
"menstruation",
"kondom",
"mens",
"mensskydd"
],
"amenity/vending_machine/food":[
"mat",
"matvarumaskin",
"matautomat",
"Matvaruautomat",
"varuautomat",
"varumaskin",
"matvaruautomat",
"mellanmål"
],
"amenity/vending_machine/fuel":[
"Bränslepump",
"diesel",
"ing",
"tanka",
"bensinstation",
"propan",
"bränslepump",
"tankomat",
"tankstation",
"mack",
"bensin",
"etanol",
"bränsle",
"tapp",
"pump",
"cng",
"biodiesel"
],
"amenity/vending_machine/ice_cream":[
"glass",
"Glassautomat",
"varuautomat",
"isglass",
"varumaskin",
"glassautomat"
],
"amenity/vending_machine/ice_cubes":[
"Ismaskin",
"varuautomat",
"is",
"varumaskin",
"iskuber",
"ismaskin"
],
"amenity/vending_machine/newspapers":[
"Tidningsautomat",
"tidning",
"tidningsdistribution",
"tidningar",
"tidningsautomat",
"tidningsutlämning",
"tidningslåda"
],
"amenity/vending_machine/parcel_pickup":[
"amazon",
"webbshop",
"paketutlämning",
"leverans",
"internetbutik",
"paketautomat",
"paketleverans",
"paket",
"utlämning",
"Paketautomat (utlämning)",
"inposts"
],
"amenity/vending_machine/parcel_pickup_dropoff":[
"amazon",
"packetinlämning",
"webbshop",
"paketutlämning",
"leverans",
"internetbutik",
"paketautomat",
"paketleverans",
"paket",
"utlämning",
"Paketautomat (ut- och inlämning)",
"inposts"
],
"amenity/vending_machine/parking_tickets":[
"parkeringsur",
"biljett",
"parkeringsavgift",
"parkeringsautomat",
"parkometer",
"parkering",
"Parkeringsautomat"
],
"amenity/vending_machine/public_transport_tickets":[
"tågbiljett",
"tågbiljetter",
"transport",
"tunnelbana",
"färja",
"båt",
"Biljettautomat för kollektivtrafik",
"bussbiljetter",
"biljett",
"biljettautomat",
"tåg",
"bussbiljett",
"spårvagn",
"buss"
],
"amenity/vending_machine/stamps":[
"porto",
"frankering",
"post",
"varuautomat",
"Frimärksautomat",
"frankeringsautomat",
"frimärksautomat",
"varumaskin",
"frimärke",
"vykort",
"brev"
],
"amenity/vending_machine/sweets":[
"tuggummi",
"tuggummiautomater",
"chips",
"godis",
"Godisautomat",
"godisautomat",
"mellanmål"
],
"amenity/veterinary":[
"veterinär",
"djurdoktor",
"djurläkare",
"djurklinik",
"djursjukhus",
"Veterinär"
],
"amenity/waste/dog_excrement":[
"hund",
"sopkärl",
"hundbajspåse",
"bajs",
"Sopkärl för hundbajspåsar",
"sopkärl för hundbajspåsar",
"hundskit",
"hundbajs",
"bajspåsar",
"skitpåse",
"hundbajspåsar",
"soptunna"
],
"amenity/waste_basket":[
"skräpkorg",
"skräp",
"Soptunna (liten)",
"sopkärl",
"papperskorg",
"papperskärl",
"avfallskorg",
"soptunna",
"sopor"
],
"amenity/waste_disposal":[
"industrisopor",
"sopkärl",
"avfall",
"avfallskärl",
"avfallstunna",
"hushållssopor",
"avfallskontainer",
"Soptunna (hushålls- eller industrisopor)",
"soptunna",
"sopor"
],
"amenity/waste_transfer_station":[
"skräp",
"avfallscentral",
"dumpa",
"skrot",
"återvinning",
"Avfallscentral"
],
"amenity/water_point":[
"dricksvatten",
"dricksvatten för campingfordon",
"vattenpåfyllning",
"Dricksvatten för campingfordon"
],
"amenity/watering_place":[
"dricksvatten",
"utfodring",
"dricksvatten för djur",
"djurutfodring",
"Dricksvatten för djur",
"vattenhåll",
"djur",
"vattenkar"
],
"amenity/weighbridge":[
"väga",
"Lastbilsvåg",
"lastbilsvåg",
"våg",
"vågstation",
"vikt",
"tyngd"
],
"area":[
"fällt",
"areal",
"område",
"utrymme",
"yta",
"Yta",
"plan",
"mark"
],
"area/highway":[
"trottoarkant",
"vägplan",
"vägbeläggning",
"Vägyta",
"vägyta",
"area:highway",
"torg",
"vägform",
"vägkant",
"köryta",
"promenatyta",
"trottoar"
],
"attraction":[
"Attraktion"
],
"attraction/amusement_ride":[
"åkattraktion",
"karusell",
"nöjespark",
"Åkattraktion",
"temapark",
"tivoli",
"nöjeskarusell"
],
"attraction/animal":[
"safari",
"Djurinhägnad",
"djurpark",
"temapark",
"fiskar",
"fågel",
"pingvin",
"tiger",
"djur",
"akvarium",
"insekt",
"djurinhägnad",
"lejon",
"djurhage",
"björn",
"apa",
"fisk",
"reptil",
"zoo",
"däggdjur",
"zoologisk trädgård"
],
"attraction/big_wheel":[
"åkattraktion",
"karusell",
"pariserhjul",
"nöjespark",
"temapark",
"stort hjul",
"tivoli",
"Pariserhjul",
"nöjeskarusell"
],
"attraction/bumper_car":[
"åkattraktion",
"Radiobilar",
"nöjespark",
"temapark",
"radiobil",
"tivoli",
"radiobilar"
],
"attraction/bungee_jumping":[
"Bungyjump",
"bungee jump",
"nöjespark",
"temapark",
"hopplattform",
"tivoli",
"bungyjump"
],
"attraction/carousel":[
"åkattraktion",
"karusell",
"nöjespark",
"temapark",
"Karusell (roterande)",
"tivoli",
"nöjeskarusell"
],
"attraction/dark_ride":[
"åkattraktion",
"karusell",
"nöjespark",
"temapark",
"tivoli",
"mörk åktur",
"spöktåg",
"nöjeskarusell",
"Mörk åktur"
],
"attraction/drop_tower":[
"fritt fall",
"åkattraktion",
"karusell",
"nöjespark",
"temapark",
"tivoli",
"nöjeskarusell",
"Fritt fall"
],
"attraction/kiddie_ride":[
"åkattraktion",
"småbarnskarusell",
"kiddie ride",
"Kiddie Ride (åkattraktion för små barn)",
"småbarnsåkattraktion"
],
"attraction/log_flume":[
"log flume",
"nöjespark",
"temapark",
"tivoli",
"stock",
"Flumeride",
"flumeride"
],
"attraction/maze":[
"slingergång",
"trojeborg",
"Labyrint",
"trojaborg",
"trädgårdslabyrint",
"labyrint",
"irrgång"
],
"attraction/pirate_ship":[
"karusell",
"nöjespark",
"temapark",
"piratskepp",
"nöjeskarusell",
"åkattraktion",
"båtgunga",
"roterande båt",
"vikingaskepp",
"gunga",
"tivoli",
"Båtgunga",
"gungande båt"
],
"attraction/river_rafting":[
"åkattraktion",
"karusell",
"nöjespark",
"forsränning",
"temapark",
"forsbana",
"fors",
"tivoli",
"Forsränning",
"vattenbana",
"nöjeskarusell"
],
"attraction/roller_coaster":[
"åkattraktion",
"berg- och dalbana",
"bergochdalbana",
"dalbana",
"Berg- och dalbana",
"nöjespark",
"temapark",
"berg-och-dalbana",
"berg-och-dal-bana",
"bergodalbana",
"tivoli"
],
"attraction/summer_toboggan":[
"kälke",
"sommerrodelbahn",
"Sommarrodel",
"rodel",
"sommarrodel",
"alpine slide",
"mountain coaster"
],
"attraction/swing_carousel":[
"åkattraktion",
"karusell",
"nöjespark",
"temapark",
"gunga",
"Gungkarusell",
"tivoli",
"gungkarusell",
"nöjeskarusell"
],
"attraction/train":[
"stadståg",
"sightseeing",
"vägtåg",
"sightseeingtåg",
"Turisttåg (ej på räls)",
"turisttåg",
"tuff tuff-tåg",
"tschu-tschu"
],
"attraction/water_slide":[
"vattenrutschkana",
"Vattenrutschbana",
"rutschkana",
"vattenrutschbana"
],
"barrier":[
"bom",
"räcke",
"avspärrning",
"stopp",
"Barriär",
"skydd",
"hinder",
"blockering",
"mur",
"barriär",
"vall",
"spärr"
],
"barrier/block":[
"trafikbarriärer",
"sugga",
"Block",
"block",
"betongsugga",
"avspärrare",
"trafikhinder"
],
"barrier/bollard":[
"stolpe",
"Stolpe",
"pollare"
],
"barrier/bollard_line":[
"stolpe",
"Stolprad",
"stolprad",
"barriär",
"pollare"
],
"barrier/border_control":[
"passkontroll",
"pass",
"tull",
"gränskontroll",
"Gränskontroll",
"säkerhetskontroll",
"gräns"
],
"barrier/cattle_grid":[
"Färist",
"färist",
"galler",
"rist"
],
"barrier/chain":[
"Kedja",
"kedja",
"kätting"
],
"barrier/city_wall":[
"skans",
"vallar",
"Stadsmur",
"befästningsverk",
"fort",
"barrikad",
"mur",
"ringmur",
"stadsmur"
],
"barrier/cycle_barrier":[
"Cykelbarriär",
"hinder",
"barriär",
"cykelbarriär"
],
"barrier/ditch":[
"dike",
"ränna",
"vallgrav",
"Dike"
],
"barrier/entrance":[
"Entré"
],
"barrier/fence":[
"gärdsgård",
"inhägnad",
"staket",
"stängsel",
"Staket"
],
"barrier/fence/railing":[
"skyddsräcke",
"trafikseparering",
"räcke",
"staket",
"Räcke",
"handräcke"
],
"barrier/gate":[
"grind",
"Grind"
],
"barrier/guard_rail":[
"kraschbarriär",
"skyddsräcke",
"krockbarriär",
"trafikseparation",
"trafikbarriär",
"kollisionsbarriär",
"Skyddsräcke"
],
"barrier/hedge":[
"Häck",
"häck",
"buskar"
],
"barrier/height_restrictor":[
"restriktion",
"höjdrestriktion",
"Höjdrestriktion",
"max",
"maxhöjd",
"höjd"
],
"barrier/kerb":[
"trottoarkant",
"kantsten",
"Trottoarkant",
"kant"
],
"barrier/kerb/flush":[
"trottoarkant",
"Trottoarkant utan upphöjning",
"trottoarkant utan upphöjning",
"kantsten",
"barnvagnsramp",
"kantstensramp",
"trottoarsramp",
"rullstolsramp",
"kant",
"nedsänkt kant",
"sluttande",
"nedsänkt trottoar",
"avfasad trottoar",
"kantstensskärning"
],
"barrier/kerb/lowered":[
"trottoarkant",
"kantsten",
"Nedsänkt trottoarkant",
"sluttande",
"nedsänkt trottoar",
"barnvagnsramp",
"kantstensramp",
"trottoarsramp",
"rullstolsramp",
"kantstensskärning",
"kant",
"nedsänkt kant"
],
"barrier/kerb/raised":[
"trottoarkant",
"upphöjd trottoar",
"kantsten",
"busshållplats",
"upphöjd kant",
"upphöjd trottoarkant",
"kant",
"Upphöjd trottoarkant"
],
"barrier/kerb/rolled":[
"trottoarkant",
"kantsten",
"Rundad trottoarkant",
"rundad trottoarkant",
"kant"
],
"barrier/kissing_gate":[
"Grind vid betesmark",
"kryssgrind",
"grind vid betesmark"
],
"barrier/lift_gate":[
"bom",
"Bom",
"avspärrning",
"lyftbom",
"spärr"
],
"barrier/retaining_wall":[
"stödmur",
"Stödmur",
"nivåskillnad"
],
"barrier/sally_port":[
"entré",
"slottsport",
"port",
"entréport",
"Befäst entréport",
"borgport",
"befäst entréport"
],
"barrier/spikes":[
"stingers",
"spikremsa",
"däckförstörare",
"Spikremsa",
"däckdeflationsanordning",
"trafikspikar",
"spikmatta",
"enkelriktning",
"stopppinnar"
],
"barrier/stile":[
"övergång",
"trappa",
"Övergång"
],
"barrier/swing_gate":[
"bom",
"Svänggrind",
"grind",
"avspärrning",
"svänggrind",
"spärr"
],
"barrier/toll_booth":[
"vägavgift",
"importavgift",
"tullmyndighet",
"gränstull",
"tullvisitation",
"tullkontroll",
"Tullstation",
"tullstation",
"tullhus",
"införselavgift",
"skatt"
],
"barrier/turnstile":[
"spärrkors",
"Vändkors",
"vändkors",
"spärr"
],
"barrier/wall":[
"befästning",
"vägg",
"hinder",
"murverk",
"mur",
"skyddsvärn",
"Mur",
"barriär"
],
"barrier/wall/noise_barrier":[
"bullerhinder",
"Ljudbarriär",
"bullerskärm",
"akustik",
"ljudhinder",
"ljudbarriär",
"buller",
"akustisk barriär",
"ljudvägg",
"akustiskt hinder",
"ljud"
],
"boundary":[
"Gräns"
],
"boundary/administrative":[
"gränslinje",
"Administrativ gräns",
"administrativ gräns",
"gräns"
],
"bridge/support":[
"pylon",
"stödpelarna",
"anfang",
"bropelare",
"landfäste",
"brostöd",
"akvedukt",
"snedkabelbro",
"Brostöd",
"stöd",
"viadukt",
"förankring",
"hängbro",
"bro"
],
"bridge/support/pier":[
"akvedukt",
"stöd",
"viadukt",
"vägport",
"överfart",
"stödpelare",
"pelare",
"balkbro",
"bro",
"Stödpelare"
],
"building":[
"anläggning",
"fastighet",
"kåk",
"byggnad",
"bygge",
"konstruktion",
"hus",
"Byggnad",
"byggnadsverk"
],
"building/apartments":[
"bostadshus",
"lägenheter",
"Lägenhetsbyggnad",
"bostad",
"lägenhetsbyggnad",
"lägenhet",
"hyreshus"
],
"building/barn":[
"lada",
"lagård",
"loge",
"ladugård",
"Lada",
"magasin",
"skjul",
"skulle"
],
"building/boathouse":[
"Båthus",
"båthus",
"sjöbod",
"strandbod"
],
"building/bungalow":[
"fristående hus",
"bungalow",
"stuga",
"sommarstuga",
"Bungalow",
"semesterhus",
"villa"
],
"building/bunker":[
"Bunker"
],
"building/cabin":[
"kåk",
"stuga",
"sommarstuga",
"Stuga",
"hus",
"koja",
"fritidshus",
"landställe",
"torp"
],
"building/carport":[
"Carport",
"garage",
"bilparkering",
"biltak",
"övertäckt parkering",
"carport",
"parkering"
],
"building/cathedral":[
"helgedom",
"dom",
"stiftskyrka",
"Katedral",
"kyrka",
"katedral",
"religiös anläggning",
"kyrkogård",
"basilika",
"kyrkobyggnad",
"religiös",
"religiöst område",
"vallfärdsort",
"gudshus",
"biskopskyrka",
"tillbedjan",
"andligt område",
"fristad",
"huvudkyrka",
"kloster",
"predikan",
"vallfärgsplats",
"kristen",
"kyrkbyggnad",
"religion",
"tro",
"kyrkorum",
"gud",
"biskop",
"dyrkan",
"guds hus",
"gudstjänst",
"kyrksal",
"domkyrka",
"kristendom"
],
"building/chapel":[
"helgedom",
"andaktssal",
"tempelområde",
"kyrka",
"religiös anläggning",
"kyrkogård",
"böneplats",
"kor",
"tempel",
"kyrkobyggnad",
"religiös",
"religiöst område",
"bönhus",
"sidokapell",
"andaktsrum",
"gudshus",
"tillbedjan",
"begravningskapell",
"fristad",
"kranskapell",
"socken",
"predikan",
"dopkapell",
"kapell",
"kristen",
"Kapell",
"kyrkbyggnad",
"mässkapell",
"religion",
"tro",
"slottskapell",
"gravkapell",
"annexkyrka",
"kyrkorum",
"mission",
"bönehus",
"andaktslokal",
"gudstjänstlokal",
"gud",
"dyrkan",
"guds hus",
"gudstjänst",
"kyrksal",
"korkapell",
"kristendom",
"missionshus",
"sanktuarium"
],
"building/church":[
"helgedom",
"församling",
"tempelområde",
"kyrka",
"katedral",
"religiös anläggning",
"kor",
"vallfärdsort",
"gudshus",
"andaktsrum",
"tillbedjan",
"begravningskapell",
"andligt område",
"fristad",
"kloster",
"dopkapell",
"kapell",
"gudstjänstslokal",
"tro",
"mission",
"bönehus",
"gud",
"dyrkan",
"guds hus",
"Kyrkobyggnad",
"kristendom",
"missionshus",
"sanktuarium",
"andaktssal",
"dom",
"kyrkogård",
"böneplats",
"basilika",
"tempel",
"kyrkobyggnad",
"religiös",
"religiöst område",
"bönhus",
"sidokapell",
"kranskapell",
"socken",
"predikan",
"vallfärgsplats",
"betel",
"kristen",
"kyrkbyggnad",
"mässkapell",
"religion",
"slottskapell",
"annexkyrka",
"gravkapell",
"kyrkorum",
"andaktslokal",
"gudstjänst",
"kyrksal",
"korkapell",
"pastorat",
"tabernakel"
],
"building/civic":[
"kommunal",
"stadshus",
"kommunhus",
"civil",
"publik",
"Kommunal byggnad",
"medborgarhus"
],
"building/college":[
"gymnasium",
"gymnasie",
"gymnasiebyggnad",
"Collegebyggnad",
"universitet"
],
"building/commercial":[
"kommersiell byggnad",
"kommersiellt",
"Kontorsbyggnad",
"affärsbyggnad",
"handelsbyggnad"
],
"building/construction":[
"byggnad under uppförande",
"bygge",
"byggnad under konstruktion",
"byggarbete",
"byggnadsplats",
"byggarbetsplats",
"byggnation",
"Byggnad under uppförande"
],
"building/cowshed":[
"kalvar",
"kostall",
"ladugård",
"ko",
"Kostall",
"mjölkstall",
"kvigor",
"tjurar",
"mjölk"
],
"building/detached":[
"enfamiljshus",
"fristående hus",
"hus",
"friliggande villa",
"Fristående hus",
"friliggande hus",
"envåningshus",
"fristående villa",
"egnahem",
"kåk",
"enbostadshus",
"småhus",
"villa"
],
"building/dormitory":[
"sovsal",
"Elevhem",
"korridorboende",
"internatskola",
"internat",
"kollektiv",
"studentkorridor",
"elevhem"
],
"building/entrance":[
"Entré/utgång"
],
"building/farm":[
"lantbruk",
"gård",
"bostadshus",
"hus",
"Mangårdsbyggnad (bostadshus på gård)",
"bostad",
"mangårdsbyggnad"
],
"building/farm_auxiliary":[
"lantbruk",
"ekonomibyggnader",
"gård",
"ladugård",
"gårdsbyggnader",
"gårdshus",
"stall",
"Gårdsbyggnader",
"lantbruksbyggnader"
],
"building/garage":[
"kallgarage",
"Garage",
"bilskjul",
"garage",
"parkeringshus",
"varmgarage",
"bilstall",
"carport"
],
"building/garages":[
"kallgarage",
"bilgarage",
"Garage",
"bilförvaring",
"bilskjul",
"parkeringshus",
"uppställningsplats",
"varmgarage",
"bilstall",
"skydd för bilar",
"carport"
],
"building/grandstand":[
"åskådarplats",
"åskådare",
"sittplats",
"Huvudläktare",
"huvudläktare",
"läktare",
"publik",
"sport"
],
"building/greenhouse":[
"vinterträdgård",
"Växthus",
"driveri",
"blomsterhus",
"orangeri",
"odlingshus",
"växthus",
"drivhus",
"växtodling"
],
"building/hangar":[
"hangar",
"flyg",
"Hangar",
"flyggarage",
"flygplan",
"hangarbyggnad"
],
"building/hospital":[
"sjukvårdsinrättning",
"klinik",
"lasarett",
"sjukhem",
"sjukstuga",
"vårdhem",
"sjukhusbyggnad",
"sjukhus",
"hospital",
"Sjukhusbyggnad",
"vårdanstalt"
],
"building/hotel":[
"hotellbyggnad",
"motell",
"hotell",
"vandrarhem",
"Hotellbyggnad",
"värdshus",
"härbärge",
"pensionat",
"gästhem"
],
"building/house":[
"enfamiljshus",
"kåk",
"bostadshus",
"enbostadshus",
"hus",
"småhus",
"Enfamiljshus",
"villa",
"parhus",
"egnahem",
"radhus"
],
"building/houseboat":[
"båt",
"hem",
"husbåt",
"Husbåt",
"bostad"
],
"building/hut":[
"barack",
"hydda",
"stuga",
"skydd",
"Koja",
"koja",
"kyffe"
],
"building/industrial":[
"lager",
"Industribyggnad",
"industribyggnad",
"industri",
"fabrik"
],
"building/kindergarten":[
"dagishus",
"förskolehus",
"kindergarten",
"förskolebyggnad",
"barnomsorg",
"dagis",
"lekskola",
"dagisbyggnad",
"daghem",
"lekis",
"förskola",
"Förskolebyggnad"
],
"building/mosque":[
"Moskébyggnad",
"islam",
"muslim",
"moskébyggnad",
"muhammedansk helgedom",
"muhammedanism",
"moské",
"minaret"
],
"building/office":[
"affärscenter",
"arbetsplats",
"Kontorsbyggnad",
"kontor",
"arbetsplatser",
"kontorsbyggnad",
"kontorsområde"
],
"building/pavilion":[
"Klubbhus",
"omklädningsrum",
"paviljong",
"klubbhus",
"idrott",
"idrottsklubb",
"sport"
],
"building/public":[
"allmän byggnad",
"publik byggnad",
"offentlig byggnad",
"Publik byggnad"
],
"building/residential":[
"flerfamiljshus",
"bostadshus",
"Bostadshus",
"boningshus",
"hyreshus"
],
"building/retail":[
"affärsbyggnad",
"detaljhandel",
"butik",
"försäljningsställe",
"Affärsbyggnad",
"varuhus",
"kiosk",
"affärshus",
"affärer"
],
"building/roof":[
"överbyggnad",
"valv",
"övertäckning",
"regnskydd",
"tak",
"Tak"
],
"building/ruins":[
"husrest",
"fornlämning",
"raserad",
"förfallen",
"ruinbyggnad",
"ödehus",
"huslämning",
"ruin",
"Ruinbyggnad"
],
"building/school":[
"gymnasium",
"skolhus",
"undervisning",
"grundskola",
"utbildning",
"skola",
"undervisningsanstalt",
"högstadium",
"folkhögskola",
"mellanstadium",
"komvux",
"skolbyggnad",
"Skolbyggnad",
"läroanstalt",
"läroverk",
"skolväsen",
"lärosäte",
"lågstadium"
],
"building/semidetached_house":[
"fristående hus",
"radhusområde",
"hus",
"friliggande hus",
"småhus",
"villa",
"parhus",
"Delvist Fristående hus",
"radhus",
"parhusområde"
],
"building/service":[
"teknikhus",
"transformator",
"nätstation",
"Teknikhus",
"teknik",
"transformatorhus",
"fördelningsstation",
"mäthus",
"pumphus",
"mätstation",
"pump",
"mätning"
],
"building/shed":[
"uthus",
"förråd",
"visthusbod",
"visthus",
"Skjul",
"förvaring",
"verkstad",
"skjul",
"förvaringsskjul",
"barack",
"hobbyhus",
"bod",
"friggebod",
"hobbyrum"
],
"building/stable":[
"stallbyggnad",
"hästar",
"ridhusanläggning",
"ridhus",
"Stall",
"stall",
"häst"
],
"building/stadium":[
"stadion",
"arenabyggnad",
"byggnad",
"friidrottsstadion",
"Stadionbyggnad",
"stadium",
"arena",
"stadionbyggnad"
],
"building/static_caravan":[
"villavagn",
"husvagn",
"campingvagn",
"Villavagn"
],
"building/sty":[
"Svinstia",
"bås",
"sugga",
"grislada",
"gris",
"svinstia",
"kulting",
"grisladugård",
"grisbås",
"svin",
"stia",
"svinladugård"
],
"building/temple":[
"fristad",
"helgedom",
"tempelområde",
"religiös anläggning",
"böneplats",
"tempel",
"religion",
"tro",
"tempelbyggnad",
"religiös",
"religiöst område",
"mission",
"Tempelbyggnad",
"bönehus",
"bönhus",
"andaktsrum",
"gudshus",
"gud",
"dyrkan",
"guds hus",
"tillbedjan"
],
"building/terrace":[
"Terrasshus",
"terrasshus"
],
"building/train_station":[
"Stationshus"
],
"building/transportation":[
"linbaneterminal",
"Byggnad för kollektivtrafik",
"färjeterminal",
"linbana",
"linjetrafik",
"terminal",
"transport",
"färja",
"båt",
"kollektivtrafikbyggnad",
"kollektivtrafik",
"bussterminal",
"båtterminal",
"spårvagnsterminal",
"metro",
"transit",
"station",
"byggnad för kollektivtrafik",
"perrong",
"buss"
],
"building/university":[
"universitetsbyggnad",
"högskola",
"Universitetsbyggnad",
"högskolebyggnad",
"universitet"
],
"building/warehouse":[
"lager",
"lada",
"lagerhus",
"upplag",
"depå",
"packhus",
"Lagerhus",
"magasin"
],
"building_part":[
"3d",
"enkla 3d-byggnader",
"Byggnadsdel",
"byggnadsdel",
"tak"
],
"building_point":[
"Byggnad"
],
"club":[
"klubblokal",
"klubb",
"föreningslokal",
"förening",
"Klubb",
"sammanslutning",
"socialt",
"sällskap"
],
"club/sport":[
"sportklubb",
"klubblokal",
"idrottsplats",
"klubb",
"idrotta",
"atlet",
"sammanslutning",
"idrottare",
"föreningslokal",
"Idrottsklubb",
"idrottsförening",
"sporta",
"förening",
"idrott",
"socialt",
"sport",
"idrottsanläggning",
"sällskap"
],
"craft":[
"hantverkare",
"hantverk",
"Hantverk",
"skrå",
"slöjd"
],
"craft/agricultural_engines":[
"jordbruksmekaniker",
"jordbruksmaskiner",
"mekaniker",
"jordbruk",
"Jordbruksmekaniker",
"skördare",
"skördetröskor",
"lantbruksmaskiner",
"traktorer",
"motormekaniker"
],
"craft/basket_maker":[
"korgslöjd",
"korgflätning",
"korgtillverkning",
"Korgtillverkare",
"korg",
"korgtillverkare"
],
"craft/beekeeper":[
"honung",
"bi",
"biodlare",
"honungstillverkning",
"biodling",
"Biodlare"
],
"craft/blacksmith":[
"konsthantverk",
"smide",
"smidesverkstad",
"smida",
"smed",
"Smed"
],
"craft/boatbuilder":[
"båtbyggeri",
"varv",
"båtbyggare",
"Båtbyggare"
],
"craft/bookbinder":[
"bokbinderi",
"bokbindning",
"bokbindare",
"bindning",
"Bokbindare",
"böcker",
"bokreparatör",
"bok"
],
"craft/brewery":[
"ölframställning",
"öl",
"Bryggeri",
"öltillverkning",
"bryggeri"
],
"craft/carpenter":[
"timmerman",
"byggnadssnickare",
"snickare",
"träarbetare",
"grovsnickare",
"Snickare"
],
"craft/carpet_layer":[
"matta",
"mattläggning",
"golv",
"mattläggare",
"golvläggare",
"Mattläggare"
],
"craft/caterer":[
"matleverantör",
"matleverans",
"catering",
"Catering",
"cateringfirma"
],
"craft/chimney_sweeper":[
"sotare",
"skorstensfejare",
"Sotare",
"rökgång",
"sotarmurre",
"skorsten"
],
"craft/cleaning":[
"flyttstäd",
"städ",
"rengöring",
"städservice",
"Städtjänst",
"städtjänst"
],
"craft/clockmaker":[
"Urmakare (väggur)",
"urmakare",
"klockmakare"
],
"craft/confectionery":[
"konfekt",
"godistillverkare",
"sötsaker",
"godisfabrik",
"choklad",
"Godistillverkare",
"godis",
"godsaker",
"konfektyrer",
"karameller",
"pastiller"
],
"craft/distillery":[
"sprittillverkning",
"mezcal",
"bourbon",
"alkohol",
"sprit",
"gin",
"destilleri",
"hembränning",
"rom",
"tequila",
"whisky",
"vodka",
"alkoholtillverkning",
"spritdryck",
"Destilleri",
"spritdestillering",
"brandy",
"alkoholdestillering",
"scotch"
],
"craft/dressmaker":[
"sömmerska",
"klädsömmare",
"Sömmerska",
"sy",
"kvinnokläder",
"klädtillverkning",
"skräddare",
"dressmaker",
"sömnad",
"klänning",
"kläder"
],
"craft/electrician":[
"systembyggare",
"kabeldragning",
"montör",
"el",
"elkraft",
"elektriker",
"elmontör",
"elreparatör",
"starkströmsmontör",
"Elektriker"
],
"craft/electronics_repair":[
"tv-service",
"tv-reparatör",
"datorreparation",
"reparation",
"skärmbyte",
"datorservice",
"telefonreparatör",
"elektronikreparation",
"reparatör",
"elektronik",
"Elektronikreparatör",
"vitvaror",
"tvättmaskinsreparatör"
],
"craft/floorer":[
"matta",
"golv",
"parkett",
"mattläggare",
"Golvläggare",
"golvläggare",
"heltäckningsmatta"
],
"craft/gardener":[
"landskapsarkitekt",
"Trädgårdsmästare",
"trädgårdsmästare",
"trädgård",
"handelsträdgård"
],
"craft/glaziery":[
"Glasmästare",
"glasblåsare",
"glas",
"fönster",
"solskydd",
"glaskonst",
"målat glas"
],
"craft/handicraft":[
"snickeri",
"hantverk",
"konsthantverk",
"textil",
"hantverksverkstad",
"Hantverksverkstad",
"hantverkare",
"vävstuga",
"handarbete",
"sömnad",
"slöjd",
"snideri",
"hemslöjd",
"vävning"
],
"craft/hvac":[
"hvac",
"ac",
"inomhusklimat",
"energiförsörjning",
"ventilation",
"sanitet",
"avlopp",
"kyla",
"vvs",
"värme",
"air condition",
"rörmokare",
"Arbetsplats för värme, ventilation och luftkonditionering",
"övervakningssystem",
"styrsystem",
"gas",
"vattenförsörjning",
"uppvärmning",
"luftkonditionering",
"tryckluft",
"vatten",
"sprinkler",
"installationsteknik"
],
"craft/insulator":[
"Isolering",
"isolering",
"ljudisolering",
"isolerare",
"värmeisolering",
"isolationsmaterial"
],
"craft/joiner":[
"finsnickare",
"snickare",
"möbler",
"träarbetare",
"slöjd",
"Finsnickare"
],
"craft/key_cutter":[
"nyckelringar",
"hänglås",
"Nyckeltillverkning",
"nyckel",
"nycklar",
"nyckelkopiering",
"nyckelring",
"nyckeltillverkning"
],
"craft/locksmith":[
"Låssmed"
],
"craft/metal_construction":[
"metallarbetare",
"Metallarbete",
"metallindustri",
"metallarbete",
"kallbearbetning",
"svets",
"svetsare",
"svetsning"
],
"craft/painter":[
"färg",
"måleriarbetare",
"Målare",
"penslar",
"tapetsering",
"måleri",
"tapetserare",
"lackering",
"målare",
"målarmästare",
"tapeter"
],
"craft/parquet_layer":[
"parkettläggare",
"golv",
"parkett",
"parkettläggning",
"golvläggare",
"Parkettläggare"
],
"craft/photographer":[
"Fotograf",
"bild",
"fotografering",
"porträttfotografering",
"bildkonst",
"porträtt",
"kamera",
"fotograf"
],
"craft/photographic_laboratory":[
"mörkrum",
"Fotoframkallning",
"kanvas",
"framkallning",
"fotoframkallning",
"foto",
"film",
"utskrift",
"filmframkallning"
],
"craft/plasterer":[
"puts",
"Putsare",
"cement",
"gips",
"väggputs",
"putsare"
],
"craft/plumber":[
"rörmontör",
"rörläggare",
"rörmokare",
"Rörmokare",
"dränering",
"vatten",
"avlopp",
"rör"
],
"craft/pottery":[
"lergods",
"krukmakare",
"Krukmakeri",
"krukgods",
"keramik",
"porslin",
"stengods",
"glasering",
"lerkärl",
"drejare",
"drejning",
"lera",
"krukmakeri",
"keramiker"
],
"craft/rigger":[
"tackling",
"rigg",
"riggare",
"segelbåt",
"segelfartyg",
"mast",
"segel",
"Riggare",
"tågvirke"
],
"craft/roofer":[
"yttertak",
"taktegel",
"takläggning",
"takpannor",
"Takläggare",
"takläggare",
"tak",
"tegel"
],
"craft/saddler":[
"läder",
"säte",
"sadelmakare",
"Sadelmakare",
"sadelmakeri",
"sadel"
],
"craft/sailmaker":[
"Segelmakare",
"segelsömnad",
"segelmakare",
"segel",
"segelmakeri"
],
"craft/sawmill":[
"Sågverk",
"trä",
"sågverk",
"virke",
"brädor",
"bräda",
"timmer",
"plank"
],
"craft/scaffolder":[
"ställningsbyggare",
"ställning",
"Ställningsbyggare",
"byggnadsställning"
],
"craft/sculptor":[
"skulptör",
"bildhuggare",
"skulpturer",
"Skulptör",
"bildsnidare",
"skulptur",
"staty"
],
"craft/shoemaker":[
"skomakare",
"skor",
"Skomakare"
],
"craft/signmaker":[
"skyltmakare",
"skyltar",
"neon",
"skylttillverkare",
"Skyltmakare",
"neonskyltar"
],
"craft/stonemason":[
"stenhuggare",
"Stenhuggare",
"stenbrott"
],
"craft/tailor":[
"Skräddare"
],
"craft/tiler":[
"plattsättare",
"plattläggare",
"golvläggare",
"Plattsättare"
],
"craft/tinsmith":[
"plåtslagare",
"tenn",
"förtennare",
"tunnplåtslagare",
"Tennsmed",
"tennsmed"
],
"craft/upholsterer":[
"möbelstoppare",
"Möbelstoppare",
"stoppning",
"tapetserare",
"möbler"
],
"craft/watchmaker":[
"Urmakare (små klockor)",
"urmakare",
"armbandsur",
"fickur",
"klockreparatör"
],
"craft/window_construction":[
"dörr",
"dörrleverantör",
"dörrar",
"glas",
"dörrinstallatör",
"fönster",
"fönstermontör",
"fönsterinstallatör",
"Fönstertillverkare",
"dörrmontör",
"fönsterleverantör",
"dörrtillverkare",
"fönstertillverkare"
],
"craft/winery":[
"vinframställnig",
"Vinfabrik",
"vineri",
"vinproduktion",
"vin",
"vinframställning",
"vinfabrik"
],
"cycleway/asl":[
"cykelbox",
"cykelstoppmarkering",
"Cykelbox",
"cykelstopp",
"asl"
],
"demolished/building":[
"Nyligen riven byggnad"
],
"disused/amenity":[
"Oanvänd facilitet"
],
"disused/railway":[
"Oanvänt järnvägsobjekt"
],
"disused/shop":[
"Nedlagd affär"
],
"embankment":[
"Vägbank"
],
"emergency":[
"Nödutrustning"
],
"emergency/ambulance_station":[
"Ambulansstation",
"räddning",
"räddningstjänst",
"ambulansstation",
"ambulans"
],
"emergency/defibrillator":[
"hjärtstartare",
"defibrillator",
"hjärthjälp",
"Defibrillator"
],
"emergency/designated":[
"Åtkomst för utryckningsfordon – Avsedd för"
],
"emergency/destination":[
"Åtkomst för utryckningsfordon – Destination"
],
"emergency/fire_alarm":[
"brandtelefon",
"Nödtelefon",
"nödtelefon"
],
"emergency/fire_extinguisher":[
"skumsläckare",
"pulversläckare",
"vattensläckare",
"vattenpost",
"eldsläckare",
"koldioxidsläckare",
"brandsläckning",
"brandpost",
"brandslang",
"Brandsläckare",
"brandsläckare",
"handbrandsläckare",
"kolsyresläckare",
"brand"
],
"emergency/fire_hose":[
"eldsläckare",
"brandsläckning",
"brandpost",
"Brandslang",
"brandslang",
"vattenpost",
"brandsläckare",
"brand"
],
"emergency/fire_hydrant":[
"brandsläckning",
"Brandpost",
"brandpost",
"vattenpost",
"brandslang"
],
"emergency/first_aid_kit":[
"brännsår",
"sårvård",
"plåster",
"sår",
"Första hjälpen",
"första hjälpen låda",
"första hjälpen kit",
"förbandslåda",
"första hjälpen",
"förband",
"bandage"
],
"emergency/landing_site":[
"nödlandningsplats",
"helikopterplatta",
"helikopter",
"helipad",
"Nödlandningsplats"
],
"emergency/life_ring":[
"livräddningsboj",
"frälsarkrans",
"Livboj",
"livräddning",
"livboj"
],
"emergency/lifeboat_station":[
"livbåt",
"Livbåtsstation",
"räddningsbåt",
"båträddning",
"livbåtsstation",
"livräddning"
],
"emergency/lifeguard":[
"Badvakt",
"cpr",
"strandvakt",
"livräddare",
"badvakt",
"lifeguard",
"räddning"
],
"emergency/mountain_rescue":[
"räddning",
"bergsräddning",
"fjällräddning",
"Fjällräddning"
],
"emergency/no":[
"Åtkomst för utryckningsfordon – Nej"
],
"emergency/official":[
"Åtkomst för utryckningsfordon – Officiellt"
],
"emergency/phone":[
"nödnummer",
"Nödtelefon",
"nödtelefon",
"alarmtelefon",
"larmtelefon",
"alarmeringscentral"
],
"emergency/private":[
"Åtkomst för utryckningsfordon – Privat"
],
"emergency/siren":[
"larm",
"siren",
"beredskapslarm",
"mistlur",
"starktonssiren",
"varning",
"flyglarm",
"Siren",
"vma",
"tyfon",
"viktigt meddelande till allmänheten",
"hesa fredrik"
],
"emergency/water_tank":[
"vattensamling",
"kris",
"reservoar",
"räddning",
"vattentorn",
"nödtank",
"brandsläckningstank",
"lagringstank",
"brandsläckning",
"vattentank för brandsläckning",
"cistern",
"tank",
"Vattentank för brandsläckning",
"brand",
"nöd",
"vatten",
"vattentank"
],
"emergency/yes":[
"Åtkomst för utryckningsfordon – Ja"
],
"entrance":[
"ingång",
"entré",
"huvudentré",
"dörr",
"utgång",
"Entré / utgång"
],
"entrance/emergency":[
"nödutgång",
"dörr",
"branddörr",
"brandutgång",
"Nödutgång",
"utgång"
],
"entrance/emergency_ward_entrance":[
"Entré till akutmottagning",
"akuten",
"akutmottagning",
"olycksmottagning",
"ambulansmottagning",
"akutavdelning",
"entré till akutmottagning"
],
"entrance/main":[
"entré",
"ingång",
"exit",
"huvudentré",
"dörr",
"Huvudentré",
"port",
"utgång",
"inträde"
],
"ford":[
"vad",
"Vadställe",
"övergångsställe",
"vadställe"
],
"ford_line":[
"Vadställe"
],
"golf/bunker":[
"bunker",
"golf",
"sandhål",
"sandfälla",
"hinder",
"Bunker",
"sandgrop"
],
"golf/cartpath":[
"golf",
"gångväg",
"gång",
"Väg för golfbil",
"golfbana",
"golfgångväg",
"stig",
"väg för golfbil",
"golfbil"
],
"golf/clubhouse":[
"golfklubb",
"Golfklubbhus",
"fritid",
"golfhus",
"kansli",
"klubbhus",
"golfkansli",
"golfklubbhus"
],
"golf/driving_range":[
"driving range",
"drivingrange",
"golf",
"driverang",
"driver",
"Driving Range",
"golfövning",
"övning"
],
"golf/fairway":[
"golf",
"fairway",
"Fairway"
],
"golf/green":[
"puttinggreen",
"golf",
"green",
"hål",
"Green"
],
"golf/hole":[
"golfhål",
"golf",
"Golfhål",
"hål"
],
"golf/lateral_water_hazard":[
"golfhinder",
"dike",
"dam",
"golf",
"vattenhinder",
"golfbana",
"sidovattenhinder",
"vattenhål",
"sjö",
"Sidovattenhinder"
],
"golf/path":[
"golf",
"gångväg på golfbana",
"gångväg",
"gång",
"golfbana",
"Gångväg på golfbana",
"golfgångväg",
"stig"
],
"golf/rough":[
"Ruff",
"ruffen",
"ruff",
"gräs"
],
"golf/tee":[
"golf",
"utslagsplats",
"tee",
"Tee"
],
"golf/water_hazard":[
"dike",
"dam",
"golf",
"vattenhinde",
"golfbana",
"Vattenhinde",
"vattenhål",
"sjö"
],
"healthcare":[
"hälsovård",
"klinik",
"institution",
"välmående",
"Hälsovård",
"doktor",
"sjukdom",
"kirurgi",
"sjuk",
"läkare",
"hälsa",
"mottagning"
],
"healthcare/alternative":[
"naturopati",
"reiki",
"tuina",
"hydroterapi",
"herbalism",
"antroposofisk",
"hypnos",
"unani",
"ayurveda",
"alternativmedicin",
"aromaterapi",
"osteopati",
"Alternativmedicin",
"shiatsu",
"tillämpad kinesiologi",
"örtmedicin",
"homeopati",
"reflexologi",
"traditionell",
"alternativ medicin",
"akupunktur"
],
"healthcare/alternative/chiropractic":[
"ryggen",
"kiropraktik",
"ryggsmärta",
"ryggrad",
"ryggbesvär",
"smärta",
"kotknackare",
"Kiropraktik (rygg)",
"kiropraktor"
],
"healthcare/audiologist":[
"audionomi",
"hörapparat",
"audionomist",
"Audionomi (hörsel)",
"öra",
"audionom",
"örat",
"hörsel",
"ljud"
],
"healthcare/birthing_center":[
"barnbördshus",
"bb",
"graviditet",
"barnafödsel",
"bäbis",
"Förlossning",
"barn",
"förlossningsavdelning",
"baby",
"förlossning",
"bebis"
],
"healthcare/blood_donation":[
"blodgivning",
"blodcentral",
"plasmaferes",
"donera blod",
"blodtransfusion",
"bloddonation",
"ge blod",
"stamcellsdonation",
"Blodgivarcentral",
"blodgivare",
"plateletpheresis",
"blodgivarcentral",
"aferes",
"blodbank"
],
"healthcare/counselling":[
"rådgivning",
"sexrådgivning",
"rådgivningscenter",
"Rådgivningscenter",
"sexualrådgivning",
"kostrådgivning"
],
"healthcare/dentist/orthodontics":[
"tandvård",
"tänder",
"Ortodontist",
"tandställning",
"tandläkare",
"tand",
"ortodontist",
"tandreglering"
],
"healthcare/hospice":[
"döende",
"död",
"hospis",
"terminalvård",
"Hospis (palliativ vård)",
"palliativ vård"
],
"healthcare/laboratory":[
"Medicinskt laboratorium",
"diagnos",
"kemi",
"blodkontroll",
"laboratoriemedicin",
"diagnosering",
"lab",
"immunologi",
"patologi",
"laboratorium",
"analys",
"medicinskt laboratorium",
"provtagning",
"genetik",
"farmakologi",
"analysrådgivning",
"mikrobiologi",
"blodanalys",
"medicinskt lab",
"transfusionsmedicin"
],
"healthcare/midwife":[
"mödrahälsovård",
"ungdomsmottagning",
"gynekolog",
"jordemo",
"ackuschörska",
"gynekologi",
"barnmorska",
"mödravårdscentra",
"Barnmorska",
"preventivmedel"
],
"healthcare/occupational_therapist":[
"ergonomi",
"terapeut",
"Arbetsterapi",
"rehabilitering",
"hjälpmedel",
"arbetsterapi",
"terapi"
],
"healthcare/optometrist":[
"korrektionsglas",
"ögon",
"glasögon",
"Optometri (ögon)",
"linser",
"syn",
"optometri",
"synhjälpmedel",
"optometrier",
"synfel",
"ögonlaser"
],
"healthcare/physiotherapist":[
"Fysioterapi (sjukgymnastik)",
"terapeut",
"fysioterapi",
"sjukgymnastik",
"fysisk",
"fysioterapeut",
"terapi"
],
"healthcare/podiatrist":[
"Podiatri (fötter)",
"fötter",
"fothälsa",
"fotkirurgi",
"naglar",
"podiatriker",
"fot",
"podiatri"
],
"healthcare/psychotherapist":[
"terapeut",
"Psykoterapi",
"psykoterapeut",
"rådgivare",
"psykolog",
"sinne",
"ångest",
"kuratorer",
"självmord",
"terapi",
"psykologisk behandling",
"mental hälsa",
"depression",
"psykoterapi"
],
"healthcare/rehabilitation":[
"Rehabilitering",
"rehab",
"terapeut",
"rehabilitering",
"terapi"
],
"healthcare/speech_therapist":[
"röst",
"språk",
"terapeut",
"Logoped (röst/tal)",
"dysfagi",
"språkstörning",
"röststörning",
"logoped",
"tal",
"terapi",
"talstörning"
],
"highway":[
"Vägobjekt"
],
"highway/bridleway":[
"rida",
"ridväg",
"ryttare",
"ridstig",
"Ridväg",
"ridning",
"häst"
],
"highway/bus_guideway":[
"spårbuss",
"guidad buss",
"Spårbuss",
"buss"
],
"highway/bus_stop":[
"Busshållplats"
],
"highway/construction":[
"stängd",
"väg avstängd",
"Avstängd väg",
"avstängd",
"väg under konstruktion",
"vägbygge",
"avstängd väg",
"vägbyggnad"
],
"highway/corridor":[
"inomhus",
"inomhuskorridor",
"korridor",
"gång",
"korridor inomhus",
"gångpassage",
"förbindelsegång",
"Korridor inomhus"
],
"highway/crossing":[
"Korsning"
],
"highway/crossing/marked":[
"övergångsställe för gående",
"vägövergång",
"vägpassage",
"gångpassage",
"Markerad gångpassage",
"markerad gångpassage",
"övergångsställe",
"gångvägspassage",
"markerat övergångsställe"
],
"highway/crossing/marked-raised":[
"vägpassage",
"markerad gångpassage",
"puckel",
"markerad gångpassage (upphöjt)",
"markerat övergångsställe",
"övergångsställe för gående",
"vägövergång",
"gångpassage",
"markerat övergångsställe (upphöjt)",
"fartpuckel",
"Markerad gångpassage (upphöjt)",
"fartgupp",
"farthinder",
"övergångsställe",
"gångvägspassage",
"gupp"
],
"highway/crossing/unmarked":[
"övergångsställe för gående",
"vägövergång",
"Omarkerad övergång",
"vägpassage",
"gångpassage",
"omarkerad gångpassage",
"övergångsställe",
"gångvägspassage",
"omarkerat övergångsställe",
"omarkerad övergång"
],
"highway/crossing/unmarked-raised":[
"vägpassage",
"omarkerat övergångsställe (upphöjt)",
"puckel",
"omarkerat övergångsställe",
"Omarkerad övergång (upphöjt)",
"omarkerad övergång (upphöjt)",
"övergångsställe för gående",
"vägövergång",
"gångpassage",
"fartpuckel",
"fartgupp",
"farthinder",
"övergångsställe",
"gångvägspassage",
"gupp",
"omarkerad övergång"
],
"highway/crossing/zebra":[
"Markerat övergångsställe"
],
"highway/crossing/zebra-raised":[
"Markerat övergångsställe (upphöjt)"
],
"highway/cycleway":[
"cykelled",
"cykelväg",
"gc-väg",
"Cykelväg",
"cykel"
],
"highway/cycleway/bicycle_foot":[
"gång- och cykelväg",
"gång och cykelväg",
"cykelväg",
"gc-väg",
"gångväg",
"gående",
"gång",
"Cykel- och gångväg",
"cykel- och gångväg",
"gångbana",
"cykelbana",
"cykel",
"cyklande",
"gcm-väg"
],
"highway/cycleway/crossing":[
"Cykelkorsning"
],
"highway/cycleway/crossing/bicycle_foot":[
"cykelväg",
"cykel- och gångkorsning",
"gång- och cykelkorsning",
"gångväg",
"gående",
"gång",
"cykelkorsning",
"gc-övergång",
"cykelpassage",
"gång och cykelkorsning",
"gångkorsning",
"gångpassage",
"cykel",
"cyklande",
"övergångsställe",
"gc-korsning",
"Cykel- och gångkorsning",
"gc-passage"
],
"highway/cycleway/crossing/marked":[
"Markerad cykelkorsning",
"cykelöverfart",
"cykelpassage",
"cykelkorsning",
"markerad cykelkorsning"
],
"highway/cycleway/crossing/unmarked":[
"cykelöverfart",
"cykelpassage",
"cykelkorsning",
"Omarkerad cykelkorsning",
"omarkerad cykelkorsning"
],
"highway/elevator":[
"hiss",
"Hiss"
],
"highway/elevator_line":[
"bergbana",
"lutning",
"Snedhiss",
"lutande hiss",
"kabelspårväg",
"vinsch",
"funikular",
"hiss",
"elevator",
"banhiss",
"lift",
"snedbanehiss",
"snedhiss"
],
"highway/emergency_bay":[
"stopp",
"uppställning",
"Nöduppställningsplats",
"nöduppställningsplats",
"haveri",
"motorstopp",
"nödtelefon",
"nödstoppplats",
"nödstopp"
],
"highway/footway":[
"gångbana",
"gångväg",
"gc-väg",
"Gångväg",
"löparbana",
"motionsspår",
"promenad"
],
"highway/footway/access_aisle":[
"åtkomstgång",
"gångväg",
"rullstolsgång",
"Åtkomstgång",
"parkeringsgång",
"lastzoon",
"handikapparkeringsåtkomstzon"
],
"highway/footway/conveying":[
"gångrullband",
"transportband för människor",
"Rullande trottoar",
"transportband",
"rullband",
"rullande gåband",
"rullande trottoar",
"rullramp",
"transportband för personer",
"rullgångbana",
"rullande gångbana",
"rulltrottoar"
],
"highway/footway/crossing":[
"Gångpassage"
],
"highway/footway/marked":[
"övergångsställe för gående",
"Markerat övergångsställe",
"vägövergång",
"vägpassage",
"gångpassage",
"markerad gångpassage",
"övergångsställe",
"gångvägspassage",
"markerat övergångsställe"
],
"highway/footway/marked-raised":[
"Markerat övergångsställe (upphöjt)",
"vägpassage",
"markerad gångpassage",
"puckel",
"markerad gångpassage (upphöjt)",
"markerat övergångsställe",
"övergångsställe för gående",
"vägövergång",
"gångpassage",
"markerat övergångsställe (upphöjt)",
"fartpuckel",
"fartgupp",
"farthinder",
"övergångsställe",
"gångvägspassage",
"gupp"
],
"highway/footway/sidewalk":[
"gångbana",
"Trottoar",
"gångväg",
"trottoar"
],
"highway/footway/unmarked":[
"övergångsställe för gående",
"vägövergång",
"Omarkerad övergång",
"vägpassage",
"gångpassage",
"omarkerad gångpassage",
"övergångsställe",
"gångvägspassage",
"omarkerat övergångsställe",
"omarkerad övergång"
],
"highway/footway/unmarked-raised":[
"vägpassage",
"omarkerat övergångsställe (upphöjt)",
"puckel",
"omarkerat övergångsställe",
"Omarkerad övergång (upphöjt)",
"omarkerad övergång (upphöjt)",
"övergångsställe för gående",
"vägövergång",
"gångpassage",
"fartpuckel",
"fartgupp",
"farthinder",
"övergångsställe",
"gångvägspassage",
"gupp",
"omarkerad övergång"
],
"highway/footway/zebra":[
"Markerat övergångsställe"
],
"highway/footway/zebra-raised":[
"Markerat övergångsställe (upphöjt)"
],
"highway/give_way":[
"utfartsregeln",
"lämna företräde",
"väjningspliktsskylt",
"utfart",
"väjningsplikt",
"Väjningsplikt",
"företräde"
],
"highway/living_street":[
"torg",
"gångfartsområde",
"Gångfartsområde",
"gårdsgata"
],
"highway/milestone":[
"milstolpe",
"postament",
"väghållningsten",
"milsten",
"Milsten"
],
"highway/mini_roundabout":[
"Minirondell",
"minirondell",
"cirkulationsplats",
"rondell",
"trafikrondell"
],
"highway/motorway":[
"motorväg",
"Motorväg",
"snabbled",
"stadsmotorväg"
],
"highway/motorway_junction":[
"motorvägspåfart",
"trafikplats",
"mot",
"avfart",
"Motorvägspåfart / -avfart",
"motorvägsavfart",
"påfart",
"vägkorsning"
],
"highway/motorway_link":[
"trafikplats",
"motorvägsanslutning",
"avfart",
"anslutning",
"påfart",
"Anslutning, motorväg"
],
"highway/passing_place":[
"mötesplats",
"passage",
"Mötesplats",
"passeringsplats",
"möte"
],
"highway/path":[
"vandring",
"gång",
"vandra",
"vandringsled",
"Stig",
"stig",
"led",
"spår",
"löparbana",
"motionsspår",
"promenad"
],
"highway/path/boardwalk":[
"gångväg",
"Spång",
"brädor",
"stig",
"plankor",
"spång",
"plankstig",
"brädväg"
],
"highway/path/informal":[
"Informell stig",
"viltstig",
"kostig",
"genväg"
],
"highway/pedestrian_area":[
"plaza",
"gångområde",
"centrum",
"gångväg",
"torg",
"gångfartsområde",
"gångfart",
"Gågateområde",
"gågata",
"gårdsgata"
],
"highway/pedestrian_line":[
"gångområde",
"affärsgata",
"centrum",
"gångväg",
"gång",
"gående",
"torg",
"gågata",
"shoppinggata",
"promenad",
"plaza",
"gångbana",
"Gågata",
"fotgängare"
],
"highway/primary":[
"primärväg",
"riksväg",
"primär väg",
"länsväg",
"Primär väg",
"huvudväg"
],
"highway/primary_link":[
"Anslutning, primär väg",
"primärväg",
"avfart",
"riksväg",
"primär väg",
"anslutning",
"påfart",
"huvudväg"
],
"highway/raceway":[
"motorracerbana",
"go-kart",
"bil*",
"f1",
"f-1",
"race*",
"formula one",
"racerbana",
"motorbana",
"gokart",
"rallybana",
"Motorracerbana",
"tävlingsbana",
"motortävling",
"rally",
"kappkörning"
],
"highway/raceway/karting":[
"go kart",
"gokart",
"motorsport",
"kartingbana",
"Kartingbana (Gokart)",
"karting",
"kart"
],
"highway/raceway/motocross":[
"motorsport",
"off-road",
"off road-bana",
"motorcross",
"off road",
"Motocrossbana",
"motorcykelbana",
"motocrossbana"
],
"highway/residential":[
"bostadsområde",
"Bostadsgata",
"gata",
"bostadsgata",
"villaväg",
"villagata"
],
"highway/rest_area":[
"rastplats",
"bensinstation",
"Rastplats"
],
"highway/road":[
"främmande",
"ospecificerad",
"Okänd väg",
"okänd väg",
"okänd",
"obekant",
"outforskad"
],
"highway/road/bridge":[
"Okänd vägbro",
"väg",
"okänd vägbro",
"bro"
],
"highway/secondary":[
"sekundär väg",
"sekundärväg",
"länsväg",
"Sekundär väg",
"huvudväg"
],
"highway/secondary_link":[
"sekundär väg",
"Anslutning, sekundär väg",
"avfart",
"sekundärväg",
"anslutning",
"länsväg",
"påfart",
"huvudväg"
],
"highway/service":[
"Serviceväg",
"bakgård",
"uppfart",
"campinggata",
"parkeringsväg",
"industriväg"
],
"highway/service/alley":[
"Gränd",
"bigata",
"gränd",
"sidogata",
"bakgata"
],
"highway/service/drive-through":[
"hämtmat",
"genomkörning",
"drive-through",
"mcdrive",
"Drive-through"
],
"highway/service/driveway":[
"uppfart",
"privat väg",
"garageinfart",
"infart",
"Uppfart",
"villaväg"
],
"highway/service/emergency_access":[
"räddningsväg",
"brandbil",
"nödväg",
"polis",
"utrymningsväg",
"utryckningsfordon",
"brandkår",
"ambulans",
"utryckningsväg",
"brandväg",
"Åtkomst för utryckningsfordon"
],
"highway/service/parking_aisle":[
"parkeringsplats",
"parkeringsväg",
"Parkeringsväg",
"parkeringsgata"
],
"highway/services":[
"rastplats",
"bensinstation",
"snabbmat",
"restaurang",
"vägmat",
"Rastplats med försäljning"
],
"highway/speed_camera":[
"fartkamera",
"fartkontroll",
"hastighetskamera",
"trafiksäkerhetskamera",
"Fartkamera"
],
"highway/steps":[
"rulltrappa",
"trappor",
"trapp",
"trappsteg",
"Trappa",
"trappa",
"trappnedgång",
"trappuppgång"
],
"highway/steps/conveying":[
"rulltrappa",
"Rulltrappa",
"trappa",
"rörlig trappa"
],
"highway/stop":[
"lämna företräde",
"stopp",
"stoppskylt",
"Stoppskylt"
],
"highway/street_lamp":[
"lyktstolpe",
"lampa",
"gatlampa",
"gatubelysning",
"belysning",
"gatuljus",
"Gatlampa"
],
"highway/tertiary":[
"sekundära länsväg",
"huvudgata",
"Tertiär väg",
"allmän väg",
"länsväg",
"tertiär väg"
],
"highway/tertiary_link":[
"huvudgata",
"Anslutning, tertiär väg",
"avfart",
"anslutning",
"länsväg",
"påfart",
"tertiär väg"
],
"highway/toll_gantry":[
"vägavgift",
"tullportal",
"vägavgiftsportal",
"portal för vägavgift",
"vägtullsportal",
"vägtull",
"portal för vägtull",
"kamera för registreringsnummer",
"portal",
"Portal för vägtull",
"automatisk vägtull"
],
"highway/track":[
"jordbruksväg",
"Jordbruks-/skogsväg",
"åkerväg",
"traktor",
"timmer",
"brandväg",
"jordbruk",
"brandgata",
"bruksväg",
"virkesväg",
"skogsmaskin",
"åker",
"traktorväg",
"skogsväg",
"timmerväg"
],
"highway/traffic_mirror":[
"trafikspegel",
"utfartspegel",
"spegel",
"hörn",
"konvex",
"Trafikspegel",
"vägspegel",
"säkerhet"
],
"highway/traffic_signals":[
"trafikljus",
"signalljus",
"Trafiksignaler",
"trafiksignal",
"ljus",
"stoppljus"
],
"highway/trailhead":[
"cykelled",
"vandring",
"ledstart",
"start av vandringsled",
"Start av led",
"led",
"vandringsstart",
"start av cykelled",
"start av led",
"spårstart"
],
"highway/trunk":[
"stamväg",
"riksväg",
"motortrafikled",
"europaväg",
"Stamväg",
"huvudväg"
],
"highway/trunk_link":[
"Anslutning, stamväg",
"avfart",
"ramp",
"anslutning",
"europaväg",
"påfart",
"huvudväg"
],
"highway/turning_circle":[
"vändplats",
"Vändplats",
"återvändsgata",
"vändplan"
],
"highway/turning_loop":[
"refug",
"Vändslinga (refug)",
"vändslinga",
"vändlop",
"vändplats"
],
"highway/unclassified":[
"mindre väg",
"oklassificerad väg",
"Mindre/oklassificerad väg",
"övrig väg",
"industrigata",
"enskild väg",
"skogsväg",
"liten väg",
"industriväg"
],
"historic":[
"historia",
"Historisk plats",
"arv",
"historik",
"historisk plats"
],
"historic/archaeological_site":[
"historia",
"utgrävning",
"Arkeologisk plats",
"ruin",
"arkeologi",
"historisk plats",
"arkeologisk plats"
],
"historic/boundary_stone":[
"gränsmärke",
"gränssten",
"Gränssten",
"milsten",
"råmärke",
"gränsröse"
],
"historic/building":[
"slott",
"historisk byggnad",
"byggnad",
"historisk",
"museum",
"sevärdighet",
"historiskt",
"Historisk byggnad"
],
"historic/castle":[
"slott",
"Slott",
"herrsäte",
"fästning",
"borg",
"palats",
"resident"
],
"historic/castle/fortress":[
"historisk fästning",
"bunker",
"befästning",
"skans",
"historisk fäste",
"fästning",
"befästningsverk",
"ringmur",
"borg",
"Historisk fästning",
"citadell",
"slott",
"försvar",
"militär",
"fortifikation",
"historiskt fort"
],
"historic/castle/palace":[
"residens",
"slott",
"kung",
"praktfull byggnad",
"kunglig bostad",
"château",
"kunglig",
"drottning",
"Palats",
"borg",
"palats",
"palä"
],
"historic/castle/stately":[
"residens",
"slott",
"Château",
"praktfull byggnad",
"château",
"slottsvin",
"adel",
"vingård",
"borg",
"palats",
"palä",
"vinslott"
],
"historic/city_gate":[
"stadsport",
"Stadsport",
"port",
"ringmur"
],
"historic/fort":[
"historisk fästning",
"bunker",
"befästning",
"skans",
"historisk fäste",
"fästning",
"befästningsverk",
"borg",
"Historiskt fort",
"citadell",
"slott",
"försvar",
"militär",
"fortifikation",
"historiskt fort"
],
"historic/manor":[
"herrskap",
"herresäte",
"Herrgård",
"adel",
"gods",
"slot",
"egendom",
"herrgård",
"mansion"
],
"historic/memorial":[
"Minnesmärke",
"monument",
"minnessten",
"minnesmärke",
"minnestavla"
],
"historic/memorial/plaque":[
"Minnestavla",
"minne",
"inskription",
"minnestavla",
"jubileumsplatta"
],
"historic/monument":[
"Monument",
"monument",
"minnesmärke"
],
"historic/pillory":[
"Historisk skampåle",
"attraktion",
"historisk skampåle",
"spöpåle",
"skampåle",
"stupa"
],
"historic/ruins":[
"husras",
"rest",
"ödehus",
"Ruiner",
"lämning",
"ruin",
"förfallen byggnad"
],
"historic/tomb":[
"grav",
"gravhög",
"Grav",
"mausoleum",
"sarkofag",
"krigsgrav",
"pyramid",
"klippgrav",
"katakomb",
"massgrav",
"krypta",
"gravvalv"
],
"historic/wayside_cross":[
"vägkors",
"kors vid väg",
"Kors vid väg",
"pilgrim",
"krucifix"
],
"historic/wayside_shrine":[
"helgedom",
"Helgedom vid väg",
"helgedom vid väg",
"pilgrim",
"helgedom längs väg"
],
"historic/wreck":[
"båt",
"vrak",
"mast",
"skrov",
"Skeppsvrak",
"skepp",
"skeppsvrak"
],
"indoor":[
"Inomhusobjekt"
],
"indoor/area":[
"inomhusområde",
"inomhus",
"område",
"Yta inomhus",
"yta",
"inomhusyta",
"yta inomhus"
],
"indoor/corridor":[
"inomhus",
"inomhuskorridor",
"korridor",
"gång",
"korridor inomhus",
"gångpassage",
"förbindelsegång",
"Korridor inomhus"
],
"indoor/corridor_line":[
"Korridor inomhus"
],
"indoor/door":[
"ingång",
"dörr",
"inomhusdörr",
"dörröppning",
"dörram",
"dörr inomhus",
"Dörr inomhus",
"utgång"
],
"indoor/elevator":[
"hiss",
"hisschakt",
"schakt",
"Innomhushisschakt",
"innomhushisschakt"
],
"indoor/room":[
"lobby",
"foajé",
"inomhusrum",
"rum",
"Rum",
"cell",
"kammare"
],
"indoor/stairs":[
"trappor",
"trapphus",
"trapp",
"steg",
"trappa",
"trappnedgång",
"inomhustrappa",
"trappuppgång",
"Inomhustrappa"
],
"indoor/wall":[
"inomhusbarriär",
"vägg",
"rumsindelning",
"rumsuppdelning",
"Vägg inomhus",
"vägg inomhus",
"barriär inomhus"
],
"internet_access/wlan":[
"Surfzon",
"wifi",
"wifi hotspot",
"wi-fi",
"hotspot",
"surfzon",
"trådlöst lokalt nät",
"wi-fi hotspot",
"öppet trådlöst nät",
"wlan",
"trådlöst nät",
"uppkopplingszon",
"fritt trådlöst nät"
],
"junction":[
"vägkorsningar",
"trafikplats",
"gatukorsning",
"Korsning",
"vägkors",
"stoppsignal",
"järnvägskorsning",
"trafiksignal",
"stoppskylt",
"korsning",
"cirkulationsplats",
"trafikkorsning",
"övergångsställe",
"rondell"
],
"landuse":[
"Markanvändning"
],
"landuse/allotments":[
"odlingslott",
"lott",
"koloniträdgård",
"kolonilott",
"koloniområde",
"Koloniområde",
"täppa"
],
"landuse/aquaculture":[
"alger",
"musselodling",
"pärlodling",
"vattenbruk",
"Akvakultur",
"akvakultur",
"skaldjur",
"fiskodling",
"vattenväxter",
"räkor",
"fisk",
"utplantering av fisk",
"ostronodling"
],
"landuse/basin":[
"Avrinningsområde"
],
"landuse/brownfield":[
"rivningstomt",
"byggtomt",
"industriområde",
"brownfield",
"rivet",
"förorenat",
"industri",
"Övergivet industriområde (Brownfield)",
"övergivet",
"ödetomt"
],
"landuse/cemetery":[
"gravfält",
"grav",
"griftegård",
"Gravfällt",
"kyrkogård",
"begravningsplats"
],
"landuse/churchyard":[
"Kyrkogård (utan gravar)"
],
"landuse/commercial":[
"shoppingområde",
"handelsområde",
"handel",
"Kommersiell område",
"kommersiellt",
"butiksområde",
"kommersiell",
"affärsområde"
],
"landuse/construction":[
"byggnad under uppförande",
"bygge",
"Byggarbetsplats",
"byggnad under konstruktion",
"byggarbete",
"byggnadsplats",
"byggarbetsplats",
"byggnation"
],
"landuse/farm":[
"Åkermark"
],
"landuse/farmland":[
"åkerfält",
"lantbruk",
"gärde",
"inäga",
"odlingsfält",
"åkerlapp",
"åkerjord",
"Åkermark",
"odling",
"fält",
"teg",
"åker",
"åkermark"
],
"landuse/farmyard":[
"lantbruk",
"gård",
"jordbruk",
"lantegendom",
"Bondgård",
"bondgård",
"lantgård"
],
"landuse/flowerbed":[
"rabatt",
"blommor",
"blomsterrabatt",
"plantering",
"Rabatt",
"blomträdgård"
],
"landuse/forest":[
"dunge",
"skogsvård",
"skogsområde",
"Skog (brukad)",
"skog",
"skogsplan",
"skogstrakt",
"träd",
"skogsdunge",
"lund",
"skogsplantering",
"timmer"
],
"landuse/garages":[
"parking",
"kallgarage",
"bilskjul",
"Garageområde",
"garage",
"varmgarage",
"garageområde",
"bilstall",
"bilplatser",
"carport"
],
"landuse/grass":[
"refug",
"mittremsa",
"Gräs",
"klippt gräs",
"gräs",
"rondell"
],
"landuse/greenfield":[
"greenfield",
"framtid",
"Planerad byggnation",
"urbanisering",
"planerad byggnation"
],
"landuse/greenhouse_horticulture":[
"vinterträdgård",
"trädgårdsodling",
"driveri",
"blomsterhus",
"orangeri",
"odlingshus",
"växthus för trädgårdsväxter",
"blomma",
"växthus",
"drivhus",
"Växthus för trädgårdsväxter",
"växtodling"
],
"landuse/harbour":[
"båt",
"kaj",
"båtterminal",
"båtplats",
"Hamn",
"hamn",
"marin"
],
"landuse/industrial":[
"industriområde",
"fabriksområde",
"Industriområde",
"fabriksdistrikt",
"industricentrum"
],
"landuse/industrial/scrap_yard":[
"metall",
"metallskräp",
"skräp",
"bil",
"fordon",
"bilskrot",
"bärgning",
"Skrotupplag",
"vrak",
"metallavfall",
"metallåtervinning",
"skrotningsanläggning",
"bildemontering",
"skrot",
"metallskrot",
"skrotupplag"
],
"landuse/industrial/slaughterhouse":[
"Slaktare",
"slakteri",
"ko",
"gris",
"fläsk",
"fjäderfän",
"slaktare",
"styckning",
"styckare",
"kalv",
"slakt",
"chark",
"styckningsanläggning",
"kyckling",
"nötkött",
"slakthus",
"kött"
],
"landuse/landfill":[
"avfallsanläggning",
"tipp",
"Soptipp",
"avskrädeshög",
"återvinningscentral",
"soptipp"
],
"landuse/meadow":[
"slåttermark",
"äng",
"Äng"
],
"landuse/orchard":[
"fruktträd",
"fruktodling",
"äppelträd",
"fruktträdgård",
"Fruktodling"
],
"landuse/plant_nursery":[
"plantskola",
"Plantskola",
"handelsträdgård"
],
"landuse/pond":[
"Damm"
],
"landuse/quarry":[
"stenbrytning",
"täkt",
"sand",
"gruva",
"utgrävning",
"sandtäckt",
"sandtag",
"sten",
"Stenbrott/Sandtag",
"stenbrott"
],
"landuse/railway":[
"banområde",
"spårväg",
"spårkorridor",
"Banområde",
"tåg",
"spårvagn",
"järnvägsområde",
"tågområde",
"tågspår",
"järnväg",
"järnvägskorridor",
"spår"
],
"landuse/recreation_ground":[
"grönområde",
"Rekreationsområde",
"parkanläggning",
"friluftsområde",
"rekreationsområde",
"parkområde",
"trädgård",
"park"
],
"landuse/religious":[
"helgedom",
"tempelområde",
"kyrka",
"religiös anläggning",
"vallfärgsplats",
"kyrkogård",
"kristen",
"Religiöst område",
"synagoga",
"böneplats",
"religion",
"tempel",
"tro",
"religiöst område",
"religiös",
"vallfärdsort",
"gud",
"dyrkan",
"tillbedjan",
"moské",
"andligt område",
"kristendom",
"moske"
],
"landuse/reservoir":[
"Reservoar"
],
"landuse/residential":[
"bostadsområde",
"lägenhetsområde",
"förort",
"villaområde",
"Bostadsområde",
"miljonområde",
"getto"
],
"landuse/residential/apartments":[
"lägenhetsområde",
"bostadsområde",
"område",
"bostadshus",
"lägenheter",
"bostad",
"lägenhet",
"hyreshus",
"lägenhetskomplex",
"Lägenhetsområde"
],
"landuse/retail":[
"försäljningsområde",
"försäljning",
"shoppingområde",
"handel",
"handelsområde",
"shoppingcenter",
"Detaljhandel",
"detaljhandel",
"affärer",
"affärsområde",
"shopping"
],
"landuse/vineyard":[
"druvor",
"château",
"vineri",
"vingård",
"vinodling",
"vin",
"vindruvor",
"vinframställning",
"vinfält",
"Vingård"
],
"landuse/winter_sports":[
"pistområde",
"skidor",
"skidområde",
"alpint",
"skidort",
"skidbacke",
"snöbrädesområde",
"vintersport",
"pist",
"skidåkning",
"vintersportområde",
"snowboardområde",
"Vintersportområde",
"snowboard"
],
"leisure":[
"Fritidsobjekt"
],
"leisure/adult_gaming_centre":[
"spelmaskiner",
"spel",
"center för vuxenspel",
"flipper",
"spelmaskin",
"vuxenspel",
"flipperspel",
"Center för vuxenspel"
],
"leisure/amusement_arcade":[
"spelhall",
"spelkonsol",
"pay-to-play-spel",
"arkadmaskin",
"flipperspel",
"arkadspel",
"Arkadhall",
"spelhus",
"arkadhall",
"arkad",
"spel",
"flipper",
"körsimulatorer",
"videospel"
],
"leisure/bandstand":[
"bandstand",
"orkester-scen",
"orkesterscen",
"paviljong",
"musikestrad",
"musikscen",
"musikpaviljong",
"estrad",
"musik",
"scen",
"Musikestrad",
"orkester"
],
"leisure/beach_resort":[
"semesteranläggning",
"turist",
"turism",
"turistanläggning",
"badort",
"Strandresort",
"rekreationsort",
"semesterresort",
"hotell",
"strand",
"kurort",
"strandresort",
"resort",
"hotellanläggning"
],
"leisure/bird_hide":[
"fågelskådargömsel",
"utsiktstorn",
"fågeltorn",
"fågelskådningstorn",
"fågelskådare",
"fågelskådning",
"fågelskådartorn",
"Torn/gömsle för fågelskådning",
"vilttorn"
],
"leisure/bleachers":[
"bänk",
"åskådarplats",
"åskådare",
"sittplats",
"Läktare",
"läktare",
"publik",
"sport"
],
"leisure/bowling_alley":[
"kägelspel",
"Bowlinghall",
"kägelsport",
"bowlinghall",
"bowling",
"bowlingbana"
],
"leisure/common":[
"fritt tillträde",
"allmänning",
"Allmänning",
"öppet område",
"allmän mark"
],
"leisure/dance":[
"rotunda",
"valls",
"foxtrot",
"folkets park",
"bal",
"salsa",
"gammaldans",
"Dansbana",
"swing",
"balsal",
"tango",
"dansbana",
"danshus",
"bugg",
"jive"
],
"leisure/dancing_school":[
"danskurs",
"foxtrot",
"vals",
"gamaldans",
"dans",
"salsa",
"swing",
"dansskola",
"tiodans",
"tango",
"dansutbildning",
"Dansskola",
"bugg",
"jive"
],
"leisure/disc_golf_course":[
"frisbeegolfbana",
"frisbee golf",
"frisbeegolf",
"Frisbeegolfbana",
"frisbee"
],
"leisure/dog_park":[
"hundpark",
"hund",
"rastgård",
"Hundpark",
"hundgård",
"kennel",
"hundrastgård"
],
"leisure/escape_game":[
"Escape Room",
"quest room",
"escape game",
"escape room",
"pusselrum",
"rymningsspel"
],
"leisure/firepit":[
"Eldstad",
"lägereld",
"eldning",
"brasa",
"eldstad",
"campingbrasa",
"lägerplats",
"eldgrop",
"grillplats",
"grill",
"grillning"
],
"leisure/fishing":[
"fiske",
"fisk",
"Fiskeplats",
"fiskeplats",
"fiskare",
"fiskevatten"
],
"leisure/fitness_centre":[
"träning",
"styrketräning",
"gym",
"fitnesscenter",
"träningslokal",
"Gym / Fitnesscenter",
"konditionsträning",
"motionsinstitut",
"styrketräningslokal"
],
"leisure/fitness_centre/yoga":[
"meditation",
"Yogastudio",
"yogastudio",
"joga",
"yoga studio"
],
"leisure/fitness_station":[
"träning",
"motion",
"fitness",
"utomhusgym",
"gym",
"naturgym",
"utegym",
"träningsbana",
"träningsspår",
"Utomhusgym"
],
"leisure/fitness_station/balance_beam":[
"träning",
"motion",
"fitness",
"Balansbom (träning)",
"balansbom",
"utomhusgym",
"gym",
"naturgym",
"utegym",
"balans"
],
"leisure/fitness_station/box":[
"hoppövning",
"träning",
"låda",
"motion",
"fitness",
"Träningsplattform/trapsteg",
"hopp",
"plattform",
"utomhusgym",
"gym",
"naturgym",
"utegym"
],
"leisure/fitness_station/horizontal_bar":[
"träning",
"pullup",
"hävräcke",
"motion",
"pull-up",
"utomhusgym",
"naturgym",
"utegym",
"räck",
"bar",
"pull up",
"Räck (träning)",
"fitness",
"gym",
"räckhäv"
],
"leisure/fitness_station/horizontal_ladder":[
"träna",
"träning",
"pullup",
"armgång",
"motion",
"stege",
"utomhusgym",
"naturgym",
"utegym",
"räck",
"pull up",
"bar",
"monkey bars",
"fitness",
"gym",
"Armgång"
],
"leisure/fitness_station/hyperextension":[
"träna",
"träning",
"motion",
"utomhusgym",
"naturgym",
"utegym",
"Ryggsträckare",
"ryggsträckare",
"rygg",
"roman chair",
"fitness",
"gym",
"rygglyft",
"hyperextension"
],
"leisure/fitness_station/parallel_bars":[
"träna",
"barr",
"träning",
"Barrpress",
"motion",
"barrpress",
"fitness",
"dips",
"utomhusgym",
"gym",
"naturgym",
"utegym"
],
"leisure/fitness_station/push-up":[
"träna",
"träning",
"push up",
"motion",
"utomhusgym",
"armhävning",
"naturgym",
"utegym",
"armhävningsstation",
"pushup",
"Armhävningsstation",
"fitness",
"gym"
],
"leisure/fitness_station/rings":[
"träna",
"träning",
"ringar",
"pullup",
"motion",
"pull-up",
"utomhusgym",
"Ringar",
"naturgym",
"utegym",
"pull up",
"fitness",
"gym"
],
"leisure/fitness_station/sign":[
"träna",
"träning",
"motion",
"fitness",
"utomhusgym",
"träningsinstruktioner",
"gym",
"instruktionsskylt",
"naturgym",
"utegym",
"skylt",
"Träningsinstruktioner"
],
"leisure/fitness_station/sit-up":[
"träna",
"crunch",
"träning",
"motion",
"sit-up-ramp. situp-ramp",
"sit up",
"utomhusgym",
"naturgym",
"utegym",
"sit-up",
"fitness",
"Situp-ramp",
"gym",
"situp"
],
"leisure/fitness_station/stairs":[
"träna",
"trappor",
"träning",
"hoppövning",
"motion",
"utomhusgym",
"naturgym",
"utegym",
"step up",
"trapp",
"steg",
"fitness",
"hopp",
"trappa",
"plattform",
"Träningstrappa",
"gym"
],
"leisure/garden":[
"odlingslott",
"örtgård",
"Trädgård",
"botanisk trädgård",
"botanik",
"plantering",
"zoologisk trädgård",
"trädgård",
"park",
"botanisk"
],
"leisure/garden/botanical":[
"botanisk trädgård",
"Botanisk trädgård",
"ovanliga växter",
"botanik",
"plantering",
"trädgård",
"botanisk",
"park",
"växtsamling"
],
"leisure/garden/community":[
"odlingslott",
"lott",
"koloniträdgård",
"kolonilott",
"koloniområde",
"Koloniområde",
"täppa"
],
"leisure/golf_course":[
"golf",
"golfcenter",
"golfbana",
"Golfbana",
"golfanläggning"
],
"leisure/hackerspace":[
"hackare",
"projekt",
"makerspace",
"hackers",
"lan",
"Hackerspace",
"hackerspace",
"hacklab"
],
"leisure/horse_riding":[
"ridskola",
"rida",
"ryttare",
"Ridskola",
"ridhus",
"ridklubb",
"ridning",
"stall",
"hästridning",
"häst",
"häst*"
],
"leisure/ice_rink":[
"hockey",
"skridsko",
"ishockeybana",
"ishockey",
"isrink",
"Skridskobana",
"ishall",
"isbana",
"skridskohall",
"skridskoåkning",
"skridskobana",
"konstisbana",
"ishockeyhall",
"curling"
],
"leisure/indoor_play":[
"bollhav",
"lekplats",
"inomhuslekland",
"Inomhuslekland",
"lekland"
],
"leisure/marina":[
"småbåt",
"båt",
"småbåtshamn",
"yacht",
"marina",
"segelbåt",
"hamn",
"fritidsbåt",
"gästhamn",
"Marina"
],
"leisure/miniature_golf":[
"minigolf",
"miniatyrgolf",
"bangolf",
"äventyrsgolf",
"Minigolf"
],
"leisure/nature_reserve":[
"reservat",
"naturpark",
"naturområde",
"nationalpark",
"Naturreservat",
"naturreservat",
"naturskyddsområde"
],
"leisure/outdoor_seating":[
"ölträdgård",
"al fresco",
"servering",
"beer garden",
"utomhusmatsal",
"restaurang",
"Uteservering",
"café",
"bar",
"utomhus",
"terrass",
"pub",
"glassbar",
"uteservering"
],
"leisure/park":[
"grönområde",
"oas",
"nöjesträdgård",
"stadsoas",
"skog",
"gräs",
"skogsmark",
"friluftsområde",
"lund",
"Park",
"plaza",
"gräsmatta",
"lekplats",
"esplanad",
"rekreationsområde",
"plantering",
"trädgård",
"park",
"äng"
],
"leisure/picnic_table":[
"bänk",
"Picknickbord",
"bord",
"matbord",
"utflyktsbord",
"picknickbord",
"picknick",
"utebord"
],
"leisure/picnic_table/chess":[
"bänk",
"shack",
"schackspelare",
"spelbord",
"schackbräda",
"schackbord",
"Schackbord"
],
"leisure/pitch":[
"stadion",
"fällt",
"idrottsplats",
"idrottsplan",
"sportplats",
"Idrottsplats",
"arena",
"plan",
"idrottsanläggning"
],
"leisure/pitch/american_football":[
"amerikansk fotbollsplan",
"amerikansk fotboll",
"football",
"Plan för amerikansk fotboll"
],
"leisure/pitch/australian_football":[
"australiensisk fotboll",
"afl",
"Australisk fotbollsplan",
"australisk fotboll",
"australisk fotbollsplan",
"aussie",
"fotboll"
],
"leisure/pitch/badminton":[
"badmintonbana",
"badminton",
"badmintonplan",
"Badmintonplan",
"fjäderboll"
],
"leisure/pitch/baseball":[
"baseballplan",
"baseball",
"Baseballplan",
"baseball-plan"
],
"leisure/pitch/basketball":[
"Basketplan",
"basket",
"basketplan",
"korgboll"
],
"leisure/pitch/beachvolleyball":[
"beachvolleyhall",
"beachfotboll",
"beachhall",
"beachvolleyplan",
"Beachvolleyplan",
"beachhandboll",
"beachvolleyboll",
"beachvolley",
"strandvolleyboll",
"volleyboll",
"beachplan"
],
"leisure/pitch/boules":[
"bocce",
"pétanque",
"boule",
"Boule/Bocce-plan",
"lyonnaise"
],
"leisure/pitch/bowls":[
"shortmat",
"bowls",
"Bowlsplan"
],
"leisure/pitch/chess":[
"schack",
"gårdsschack",
"Stort schackbräde",
"schackbräde",
"parkschack",
"stort schackbräde",
"schackbord",
"schackbräda",
"trädgårdsschack"
],
"leisure/pitch/cricket":[
"kricket",
"cricket",
"Cricketplan",
"cricketplan",
"kricketplan"
],
"leisure/pitch/equestrian":[
"ridskola",
"rida",
"trav",
"ridhus",
"ridklubb",
"Ridområde",
"ridning",
"stall",
"dressyr",
"häst",
"häst*",
"galopp",
"ryttare",
"hästridning",
"hästhoppning"
],
"leisure/pitch/field_hockey":[
"landhockey",
"Landhockeyplan",
"landhockeyplan"
],
"leisure/pitch/horseshoes":[
"Kasta hästsko",
"kasta hästsko",
"hästsko"
],
"leisure/pitch/netball":[
"Nätbollsplan",
"basket",
"nätbollsplan",
"nätboll",
"dambasket",
"netball"
],
"leisure/pitch/rugby_league":[
"rugby football",
"rugby",
"rugger",
"rugbyplan",
"rugby league",
"Rugby League-plan"
],
"leisure/pitch/rugby_union":[
"Rugby Union-plan",
"rugby football",
"rugby union-plan",
"rugby",
"rugger",
"rugbyplan",
"rugby union"
],
"leisure/pitch/shuffleboard":[
"golvshuffleboard",
"bordsshuffleboard",
"Shuffleboardbana",
"shuffleboard",
"shuffleboardbana"
],
"leisure/pitch/skateboard":[
"skateboardramp",
"halfpipe",
"skateboard",
"Skateboardpark",
"skateboardpark",
"skate park"
],
"leisure/pitch/soccer":[
"fotbollsplan",
"Fotbollsplan",
"fotboll"
],
"leisure/pitch/softball":[
"softball",
"baseboll",
"brännboll",
"Softballplan",
"softballplan",
"boboll"
],
"leisure/pitch/table_tennis":[
"ping pong",
"bordtennisbord",
"pingis",
"bordtennis",
"pingpongbord",
"Pingisbord",
"pingpong",
"pingisbord"
],
"leisure/pitch/tennis":[
"tennisbana",
"Tennisbana",
"tennis",
"tennisplan"
],
"leisure/pitch/volleyball":[
"volleybollplan",
"beachvolleyboll",
"Volleybollplan",
"volleyboll"
],
"leisure/playground":[
"Lekplats",
"lek",
"lekplats",
"lekområde",
"klätterställning",
"gunga",
"lekpark"
],
"leisure/playground/indoor":[
"bollhav",
"lekplats",
"Inomhuslekplats",
"inomhuslekplats",
"lekland"
],
"leisure/resort":[
"semesteranläggning",
"rekreationsort",
"turist",
"semesterresort",
"hotell",
"Resort",
"kurort",
"turism",
"turistanläggning",
"resort",
"badort",
"hotellanläggning"
],
"leisure/sauna":[
"kölna",
"badstuga",
"bastu",
"sauna",
"Bastu"
],
"leisure/slipway":[
"sjösättning",
"Stapelbädd",
"båtramp",
"staplar",
"sjösättningsplats",
"varv",
"docka",
"torrdocka",
"stapelbädd",
"fartygsdocka"
],
"leisure/slipway_point":[
"sjösättning",
"båtramp",
"Sjösättningsplats",
"staplar",
"sjösättningsplats",
"varv",
"docka",
"torrdocka",
"stapelbädd",
"fartygsdocka"
],
"leisure/sports_centre":[
"idrottsplats",
"träning",
"sportanläggning",
"idrottsplan",
"motion",
"träningsanläggning",
"fitnes",
"sportpalats",
"idrottshall",
"Sportcenter / -anläggning",
"gym",
"simhall",
"sportcenter",
"sporthall",
"idrottsanläggning"
],
"leisure/sports_centre/climbing":[
"firning",
"klättringsgym",
"klättring",
"repellering",
"klättervägg",
"bouldering",
"bergsvägg",
"topprepsklättring",
"klättergym",
"repklättring",
"Klättergym",
"konstgjord klättervägg",
"topprep",
"rep",
"bergsklättring"
],
"leisure/sports_centre/swimming":[
"badhus",
"simbassäng",
"badhall",
"simning",
"pool",
"tävlingssim",
"Badanläggning",
"badanläggning",
"simhall",
"bassäng",
"swimmingpool",
"motionssim"
],
"leisure/sports_hall":[
"inomhusidrott",
"sportarena",
"idrottshall",
"gym",
"sporthall",
"Sporthall"
],
"leisure/stadium":[
"Stadium",
"stadium",
"arena"
],
"leisure/swimming_area":[
"naturbad",
"strand",
"badstrand",
"bad",
"dyka",
"naturbadområde",
"klippbad",
"badsjö",
"vatten",
"Naturbadområde"
],
"leisure/swimming_pool":[
"Simbassäng",
"simbassäng",
"simning",
"pool",
"bassäng",
"swimmingpool",
"simma"
],
"leisure/track":[
"cykeltävling",
"cykellopp",
"kapplöpningsbana",
"travbana",
"Tävlingsbana (Icke motorsport)",
"hundkapplöpning",
"löpbana",
"galoppbana",
"tävlingsbana",
"hästkapplöpning",
"löpning"
],
"leisure/track/cycling":[
"cykelväg",
"cykelspår",
"cykel",
"cykelbana",
"Tävlingsbana (Cykel)",
"cykelstig"
],
"leisure/track/horse_racing":[
"kapplöpning",
"galopp",
"kapplöpningsbana",
"trav",
"Tävlingsbana (Hästkapplöpning)",
"hästkapplöpningsbana",
"hästkapplöpning",
"häst"
],
"leisure/track/running":[
"kapplöpningsbana",
"sprint",
"språng",
"springa",
"Tävlingsbana (Löpning)",
"löpbana",
"tävlingsbana",
"löpning",
"löparbana"
],
"leisure/trampoline_park":[
"hoppa",
"trampolinpark",
"studsa",
"Trampolinpark",
"studsmatta",
"trampolin"
],
"leisure/water_park":[
"vattenpark",
"vattenland",
"Äventyrsbad / Vattenpark",
"äventyrsbad",
"vattenlekpark"
],
"line":[
"utsträckning",
"sträcka",
"streck",
"Linje",
"linje"
],
"man_made":[
"Människoskapat objekt"
],
"man_made/adit":[
"gruvhål",
"gruvingång",
"stoll",
"gruva",
"gruvgång",
"horisontell gruvgång",
"Horisontell gruvgång (Stoll)",
"stollen",
"lichtloch",
"dagort",
"sidoort"
],
"man_made/antenna":[
"mobil",
"Antenn",
"mobilmast",
"tv",
"antenn",
"överföring",
"mast",
"sändning",
"radiomast",
"tv-mast",
"kommunikation",
"radio"
],
"man_made/beacon":[
"vårdkase",
"beacon",
"fyrbåk",
"böte",
"Fyrbåk",
"båk",
"sjömärke",
"ledfyr",
"fyr"
],
"man_made/beehive":[
"honung",
"bikupa",
"bi",
"pollinisation",
"Bikupa",
"pollinering",
"bifarm"
],
"man_made/breakwater":[
"fördämning",
"hamnarm",
"vågbrytare",
"Vågbrytare",
"pir",
"vågskydd",
"hamnpir"
],
"man_made/bridge":[
"vägport",
"förbindelse",
"spång",
"fällbro",
"broyta",
"akvedukt",
"övergång",
"vridbro",
"viadukt",
"överfart",
"broområde",
"Broyta",
"bro"
],
"man_made/bunker_silo":[
"lager",
"spannmålssilo",
"spannmål",
"ensilage",
"pressfoder",
"foder",
"fodersilo",
"Plansilo",
"plansilo",
"silo",
"djurfoder",
"spannmålslagring"
],
"man_made/cairn":[
"röse",
"råmärken stenar",
"stenstapel",
"Stenröse",
"stenrös",
"röjningsröse",
"stenröse",
"stenhög",
"rös",
"gränsrösen"
],
"man_made/chimney":[
"Skorsten",
"rökgång",
"skorsten"
],
"man_made/clearcut":[
"föryngringsavverkning",
"skog",
"hygge",
"trä",
"träd",
"kalhygge",
"Kalhygge",
"timmer",
"avverkning",
"föryngringsyta",
"avskogning",
"slutavverkning",
"skövlat skogsområde",
"avverkningsområde"
],
"man_made/courtyard":[
"gård",
"Innergård",
"innergård",
"gårdsplan",
"torg",
"borggård",
"innetorg",
"inhägnad öppet område"
],
"man_made/crane":[
"kran",
"Kran",
"vinsch",
"travers",
"lyftkran",
"telfer"
],
"man_made/cross":[
"vägkors",
"Kors",
"kors",
"kristet kors",
"pilgrim",
"jesuskors",
"krucifix",
"kristendom"
],
"man_made/cutline":[
"pipelinegata",
"jaktgata",
"skiljelinje",
"skogssektion",
"Snittlinje i skog",
"pipeline",
"rörgata",
"gränslinje",
"skogsområde",
"brandgata",
"snittlinje",
"skidspår",
"domän",
"gräns",
"rågång"
],
"man_made/dovecote":[
"duvor",
"duva",
"brevduvor",
"duvbostad",
"Duvslag",
"fågel",
"fågelholk",
"fåglar",
"duvhus",
"duvslag"
],
"man_made/dyke":[
"fördämningsvall",
"flodvall. vattenvall",
"skyddsvall",
"vall",
"Vall (mot vatten)",
"strandvall"
],
"man_made/embankment":[
"bank",
"upphöjning",
"Vägbank",
"barnvall",
"vall",
"vägbank"
],
"man_made/flagpole":[
"Flaggstång",
"flaggstång",
"flagga"
],
"man_made/gasometer":[
"gasbehållare",
"Gasklocka",
"gasometer",
"gascistern",
"gasklocka",
"gas",
"cistern",
"stadsgas",
"naturgas"
],
"man_made/goods_conveyor":[
"Transportband",
"transportband",
"transportörsystem",
"bandtransportörer och palltransportörsystem",
"rullbanor"
],
"man_made/groyne":[
"Hövd, vågbrytare vinkelrätt mot kusten",
"vågbrytare",
"pir",
"erosion",
"hövd",
"erosionsskydd"
],
"man_made/lighthouse":[
"fyrtorn",
"fyrskepp",
"fyr",
"Fyr"
],
"man_made/manhole":[
"gatubrunn",
"dagvatten",
"telefoni",
"dagvattenbrunn",
"manhålslucka",
"Gatubrunn",
"manlucka",
"avlopp",
"telekom",
"brunnslock",
"a-brunn",
"brandpost",
"rensbrunn",
"avloppsbrunn",
"brunn",
"manhål"
],
"man_made/manhole/drain":[
"Dagvattenbrunn",
"dagvatten",
"dagvattenbrunn",
"avrinning",
"regnvatten",
"brunn",
"regn",
"avlopp"
],
"man_made/manhole/gas":[
"manhålslucka för gas",
"brunnslock",
"gatubrunn",
"gas",
"manhålslucka",
"gas-brunn",
"manlucka",
"Gatubrunn för gas",
"brunn",
"manhål"
],
"man_made/manhole/power":[
"brunnslock",
"el-brunn",
"ström",
"Manhålslucka för elkraft",
"gatubrunn",
"manhålslucka för elkraft",
"el",
"elkraft",
"manhålslucka",
"manlucka",
"brunn",
"manhål"
],
"man_made/manhole/sewer":[
"brunnslock",
"manhålslucka för avlopp",
"gatubrunn",
"manhålslucka",
"Manhålslucka för avlopp",
"manlucka",
"avloppsbrunn",
"brunn",
"avlopp",
"manhål"
],
"man_made/manhole/telecom":[
"kabel",
"manhålslucka för telekom",
"gatubrunn",
"telekom-brunn",
"telefoni",
"manhålslucka",
"manlucka",
"telekabel",
"telekom",
"brunnslock",
"telefon",
"Manhålslucka för telekom",
"tele",
"brunn",
"manhål"
],
"man_made/manhole/water":[
"dricksvatten",
"brunnslock",
"manhålslucka för vattenförsörjning",
"gatubrunn",
"vatenbrunn",
"manhålslucka",
"vattenförsörjning",
"manlucka",
"vatten",
"Manhålslucka för vattenförsörjning",
"brunn",
"manhål"
],
"man_made/mast":[
"mobiltelefon torn",
"mobilmast",
"stagas torn",
"överföringsmast",
"antennbärare",
"mast",
"mobiltelefonmast",
"radiomast",
"sändarmast",
"Mast",
"antenn",
"sändarstation",
"slavsändare",
"kommunikationsmast",
"tv-mast",
"tv-torn",
"kommunikationstorn",
"överföringstorn"
],
"man_made/mast/communication":[
"mobilmast",
"överföringsmast",
"radiomast",
"mast",
"radiotorn",
"sändartorn",
"mobilantenn",
"mobiltelefon",
"radiosändning",
"antenn",
"kommunikationsmast",
"transmissionsmast",
"radioantenn",
"Kommunikationsmast",
"tv-mast",
"tv-torn",
"kommunikationstorn",
"överföringstorn"
],
"man_made/mast/communication/mobile_phone":[
"mobilantenn",
"mobiltelefon",
"mobilmast",
"antenn",
"överföringsmast",
"Mobilmast",
"kommunikationsmast",
"transmissionsmast",
"mast",
"kommunikationstorn",
"överföringstorn"
],
"man_made/mast/communication/radio":[
"radiosändning",
"antenn",
"överföringsmast",
"transmissionsmast",
"radiomast",
"mast",
"radiotorn",
"Radiomast",
"radioantenn",
"sändartorn",
"överföringstorn"
],
"man_made/mast/communication/television":[
"mobilmast",
"tv",
"överföringsmast",
"mast",
"radiomast",
"television",
"tv-sändning",
"sändartorn",
"mobilantenn",
"mobiltelefon",
"antenn",
"kommunikationsmast",
"transmissionsmast",
"radioantenn",
"TV-mast",
"tv-mast",
"tv-torn",
"kommunikationstorn",
"överföringstorn"
],
"man_made/mineshaft":[
"grotta",
"gruvschakt",
"gruva",
"gruvgång",
"underjordisk",
"tunnel",
"Gruvschakt"
],
"man_made/monitoring_station":[
"vattennivå",
"radon",
"väderstation",
"trafik",
"väder",
"luftkvalitet",
"observation",
"övervakningsstation",
"observationsrör",
"luftkvalité",
"Mätstation",
"gps",
"jordbävning",
"trafikmätning",
"seismolog",
"seismologi",
"mätstation",
"luftmätning",
"mätning",
"ljud"
],
"man_made/obelisk":[
"obelisk",
"pelare",
"Obelisk"
],
"man_made/observatory":[
"astronomisk",
"astronom",
"meteorologisk",
"Observatorium",
"observatorium",
"rymd",
"teleskop"
],
"man_made/petroleum_well":[
"olja",
"oljetorn",
"oljeborr",
"Oljeborr",
"oljepump",
"petroleum",
"oljeborrning"
],
"man_made/pier":[
"hamnarm",
"vågbrytare",
"kaj",
"pir",
"Pir",
"hamnpir"
],
"man_made/pier/floating":[
"brygga",
"Flytande pir",
"hamnarm",
"strandpromenad",
"vågbrytare",
"kaj",
"flytande pir",
"pir",
"flytande brygga",
"hamnpir"
],
"man_made/pipeline":[
"pipeline",
"ledning",
"oljeledning",
"avloppsledning",
"vattenledning",
"rörledning",
"Pipeline"
],
"man_made/pipeline/underground":[
"olja",
"avloppsrör",
"oljepipeline",
"underjordiskt rör",
"underjordisk pipeline",
"Underjordisk pipeline",
"naturgas",
"rör",
"avlopp",
"pipeline",
"gas",
"vatten",
"vattenrör"
],
"man_made/pipeline/valve":[
"olja",
"pipelineventil",
"kran till pipeline",
"kran",
"ventil",
"kran till rör",
"gas",
"Kran till pipeline",
"pipelinekran",
"naturgas",
"vatten",
"avlopp"
],
"man_made/pumping_station":[
"vattenpump",
"avloppspump",
"Pumpstation",
"oljepump",
"spillvattenspump",
"pump",
"pumpstation",
"dräneringspump",
"pumpaggregat"
],
"man_made/reservoir_covered":[
"övertäckt reservoar",
"vattenreservoar",
"underjordisk reservoar",
"Övertäckt reservoir",
"vattentank"
],
"man_made/silo":[
"lager",
"spannmålssilo",
"spannmål",
"ensilage",
"pressfoder",
"foder",
"fodersilo",
"silo",
"Silo",
"djurfoder",
"spannmålslagring"
],
"man_made/storage_tank":[
"reservoar",
"vattentorn",
"cistern",
"Lagringstank",
"tank",
"lagringstank"
],
"man_made/storage_tank/water":[
"vattencistern",
"vattenlager",
"cistern",
"vattentorn",
"Vattentank",
"vattentank"
],
"man_made/street_cabinet":[
"gatuskåp",
"kabeltv",
"teknikskåp",
"kopplingsskåp",
"teleskåp",
"Teknikskåp",
"trafikljuskontroll",
"telefoni",
"övervakning",
"kabel-tv",
"elskåp",
"telekommunikation"
],
"man_made/surveillance":[
"övervakningsutrustning",
"bevakningskamera",
"övervakning",
"bevakning",
"övervakningskamera",
"kamera",
"Övervakning"
],
"man_made/surveillance/camera":[
"alpr",
"registreringsskylt",
"anpr",
"webbkamera",
"vakt",
"övervakning",
"Övervakningskamera",
"video",
"cctv",
"kamera",
"webcam säkerhetskamera",
"säkerhet"
],
"man_made/survey_point":[
"fixpunkt",
"Trianguleringspunkt",
"triangulering",
"trianguleringspunkt",
"kartritning"
],
"man_made/torii":[
"torii",
"jinja",
"japansk port",
"Torii",
"shinto shrine",
"fågelsittpinne",
"shintohelgedom"
],
"man_made/tower":[
"Torn",
"torn",
"radiotorn"
],
"man_made/tower/bell_tower":[
"klockgavel",
"Klocktorn",
"kyrkklocka",
"klockstapel",
"klocktorn",
"kampanil",
"kyrktorn",
"klockspel"
],
"man_made/tower/communication":[
"mobilmast",
"överföringsmast",
"radiomast",
"mast",
"radiotorn",
"sändartorn",
"mobilantenn",
"mobiltelefon",
"radiosändning",
"antenn",
"kommunikationsmast",
"transmissionsmast",
"radioantenn",
"tv-mast",
"Kommunikationstorn",
"tv-torn",
"kommunikationstorn",
"överföringstorn"
],
"man_made/tower/cooling":[
"elkraftverk",
"kolkraftverk",
"Kyltorn",
"kraftverk",
"kyltorn",
"kraftstation",
"elkraftstation",
"kärnkraftverk"
],
"man_made/tower/defensive":[
"torn",
"befästning",
"försvar",
"borgtorn",
"befästningstorn",
"befäst torn",
"försvarstorn",
"borg",
"Befäst torn"
],
"man_made/tower/minaret":[
"minâra",
"islam",
"muslim",
"böneutropare",
"muezzin",
"bönetorn",
"Minaret",
"moské",
"muaddhin",
"minaret"
],
"man_made/tower/observation":[
"utsiktstorn",
"observationstorn",
"utsiktspost",
"utkikstorn",
"observationspost",
"Utkikstorn",
"brandtorn"
],
"man_made/tower/pagoda":[
"kinesiska pagoder",
"tempeltorn",
"buddhistisk tempelbyggnad",
"buddistiskt torn",
"asiatiskt tempel",
"gudstjänstbyggnad",
"stupor",
"pagod",
"stupa",
"Pagod",
"tempel"
],
"man_made/tunnel":[
"underpassage",
"Tunnelområde",
"tunnelområde",
"underjordisk passage",
"underjordisk",
"tunnel"
],
"man_made/utility_pole":[
"elstolpe",
"elledningsstolpe",
"stolpe",
"El-/Telefonstolpe",
"telefonstolpe",
"kraftledningsstolpe"
],
"man_made/wastewater_plant":[
"avloppsreningsverk",
"reningsverk",
"avloppsverk",
"vattenreningsverk",
"Avloppsreningsverk",
"vattenrening",
"avlopp"
],
"man_made/water_tap":[
"dricksvatten",
"vattenkälla",
"vattenkran",
"kran",
"Vattenkran",
"vattenfontän",
"vattenpunkt",
"vatten"
],
"man_made/water_tower":[
"vattenreservoar",
"Vattentorn",
"vattentorn",
"vatten"
],
"man_made/water_well":[
"Brunn",
"källa",
"vattenbrunn",
"grundvatten",
"vattenhål",
"brunn"
],
"man_made/water_works":[
"vattenreningsanläggning",
"vattenreningsverk",
"vatten",
"vattenverk",
"vattenanläggning",
"Vattenverk"
],
"man_made/watermill":[
"vattenkvarn",
"vattenmölla",
"kvarnhjul",
"kvarn",
"mölla",
"skovelhjul",
"skvalta",
"Vattenkvarn",
"skvaltkvarn"
],
"man_made/windmill":[
"Väderkvarn",
"väderkvarn",
"vindmölla",
"kvarn",
"mölla",
"vädemölle",
"vindkraft"
],
"man_made/windpump":[
"vindpump",
"vattenpump",
"väderkvarn",
"aerorotor",
"vindkraftverk",
"pump",
"vindkraft",
"vind",
"Vindpump"
],
"man_made/works":[
"fabriksbyggnad",
"bil",
"bearbetningsanläggning",
"montering",
"monteringsanläggning",
"fabrikstillverkning",
"verkstad",
"raffinaderi",
"Fabrik",
"oljeraffinaderi",
"tillverkning",
"plast",
"industri",
"möbeltillverkning",
"bryggeri",
"bearbetning",
"fabrik"
],
"marker":[
"platta",
"post",
"markör",
"milsten",
"stolpe",
"märkning",
"Markör",
"identifierare",
"skylt"
],
"marker/utility":[
"platta",
"markör",
"markör av samhällsservice",
"oljeledning",
"stolpe",
"märkning",
"markör av gasledning",
"Markör av samhällsservice",
"skylt",
"rörmarkering",
"post",
"oljemarkör",
"ledningsmarkering",
"gas",
"ledningsmarkör",
"identifierare",
"markör av oljeledning"
],
"marker/utility/power":[
"platta",
"markör",
"stolpe",
"märkning",
"Kraftledningsmarkör",
"skylt",
"markör av kraftledning",
"kraftledning",
"markering av kraftledning",
"post",
"elledning",
"identifierare",
"kraftledningsmarkör"
],
"natural":[
"Naturobjekt"
],
"natural/bare_rock":[
"Kala klippor",
"klippor",
"berghäll",
"häll",
"kala klippor"
],
"natural/bay":[
"bukt",
"vik",
"Vik"
],
"natural/beach":[
"strandlinje",
"strand",
"badstrand",
"flodstrand",
"sandstrand",
"badställe",
"Strand",
"grusstrand",
"badplats"
],
"natural/cape":[
"bukt",
"udde",
"Kap (stor udde)",
"erosion",
"vik",
"kust",
"kap",
"cape"
],
"natural/cave_entrance":[
"grotta",
"bergrum",
"berghåla",
"bergsöppning",
"Grottingång",
"grotthål",
"grottöppning",
"grottingång",
"grottsystem"
],
"natural/cliff":[
"klippa",
"klippavsats",
"Klippa",
"terrass",
"stup",
"platå",
"brant",
"bergskam"
],
"natural/coastline":[
"strand",
"kustlinje",
"kustremsa",
"ö",
"kust",
"Kustlinje",
"hav"
],
"natural/fell":[
"fjäll",
"fjällandskap",
"trädgräns",
"högfjäll",
"Fjäll"
],
"natural/geyser":[
"gejser",
"het källa",
"varmvatten",
"källa",
"ånga",
"hydrogeologi",
"Gejser",
"hydrotermisk explosion"
],
"natural/glacier":[
"landis",
"jökel",
"glaciär",
"gletscher",
"ismassa",
"Glaciär"
],
"natural/grassland":[
"grässlätt",
"Grässlätt",
"gräsfällt",
"äng"
],
"natural/heath":[
"tundra",
"slätt",
"alvar",
"hed",
"kalmark",
"Hed",
"slättmark",
"gräs",
"äng",
"stäpp"
],
"natural/hot_spring":[
"gejser",
"het källa",
"termalkälla",
"Het källa"
],
"natural/mud":[
"sörja",
"sankmark och sumpmark",
"dy",
"våtmark",
"gegga",
"lera",
"gyttja",
"Lera",
"lerigt"
],
"natural/peak":[
"kulle",
"höjdpunkt",
"alp",
"hjässa",
"bergstopp",
"topp",
"berg",
"klint",
"kalott",
"Bergstopp",
"höjd",
"klätt",
"klack"
],
"natural/reef":[
"grund",
"rev",
"Rev",
"sandbank",
"undervattensgrund",
"sandrev",
"sand",
"undervattensskär",
"bank",
"korall",
"barriär",
"hav",
"revel",
"korallrev"
],
"natural/ridge":[
"kulle",
"horst",
"kam",
"berg",
"höjd",
"högland",
"bergsområde",
"krön",
"ås",
"bergsrygg",
"Ås"
],
"natural/rock":[
"klippa",
"klippa/stenbumling fäst i berggrund",
"stenbumling",
"berggrund",
"sten",
"bumling",
"Klippa/stenbumling fäst i berggrund"
],
"natural/saddle":[
"Bergskam",
"bergskrön",
"berg",
"bergskam",
"dal",
"dalgång"
],
"natural/sand":[
"sand",
"strand",
"Sand",
"öken"
],
"natural/scree":[
"stensamling",
"röse",
"lösa block",
"stenanhopning",
"Stensamling",
"block",
"taluskon",
"stenras"
],
"natural/scrub":[
"busksnår",
"sly",
"buskskog",
"snår"
],
"natural/shingle":[
"klapperstensfält",
"strand",
"klappersten",
"småsten",
"Grus (singel)",
"grus",
"rundade stenfragment",
"singel",
"flodbädd"
],
"natural/shrub":[
"Buskmark",
"buskage",
"buskmark",
"buskar"
],
"natural/spring":[
"källsprång",
"springflöde",
"Källa",
"källåder",
"källa",
"vattenställe",
"källdrag",
"källflöde",
"vattenhål"
],
"natural/stone":[
"klippa",
"klippa/stenbumling friliggande",
"friliggande sten",
"stenbumling",
"sten",
"Klippa/stenbumling friliggande"
],
"natural/tree":[
"lövträd",
"ek",
"trä",
"träd",
"barrträd",
"gran",
"Träd",
"stam",
"stock",
"trädstam",
"björk"
],
"natural/tree_row":[
"trädrad",
"boulevard",
"allé",
"aveny",
"trädkantad väg",
"Trädrad",
"lövgång",
"träallé",
"esplanad"
],
"natural/valley":[
"dal",
"sänka",
"Dal",
"dalgång"
],
"natural/volcano":[
"lava",
"vulkan",
"berg",
"vulkankrater",
"magma",
"krater",
"Vulkan"
],
"natural/water":[
"vattensamling",
"damm",
"reservoar",
"Vatten",
"göl",
"tjärn",
"vatten",
"sjö"
],
"natural/water/basin":[
"infiltrering",
"dagvatten",
"bassäng",
"Avrinningsområde",
"avrinning",
"dagvattenbassäng",
"avrinningsområde",
"infiltration"
],
"natural/water/canal":[
"vattenväg",
"ränna",
"kanal",
"vattenled",
"vattendrag",
"kanalområde",
"segelränna",
"å",
"Kanalområde",
"farled"
],
"natural/water/lake":[
"insjö",
"vattensamling",
"lagun",
"pöl",
"tjärn",
"göl",
"vatten",
"sjö",
"Sjö",
"innanhav"
],
"natural/water/moat":[
"kanal",
"Vallgrav",
"vallgrav"
],
"natural/water/pond":[
"damm",
"kvarndamm",
"Tjärn",
"liten sjö",
"tjärn",
"göl"
],
"natural/water/reservoir":[
"fördämning",
"Reservoar",
"damm",
"reservoar",
"tank"
],
"natural/water/river":[
"vattendrag",
"vattenled",
"ström",
"jokk",
"å",
"flodområde",
"fors",
"flod",
"Flodområde",
"älv"
],
"natural/water/stream":[
"dike",
"biflod",
"vattendrag",
"flöde",
"ström",
"bäck",
"biflöde",
"flod",
"bäckområde",
"rännil",
"Bäckområde"
],
"natural/water/wastewater":[
"reningsverk",
"skit",
"Avloppsvattenbassäng",
"reningsbassäng",
"avföring",
"avloppsvatten",
"avloppsvattenbassäng",
"segmenteringsbassäng"
],
"natural/wetland":[
"mad",
"Våtmark",
"sump",
"moras",
"sankmark",
"myr",
"mosse",
"träsk",
"våtmark",
"torvmark",
"kärr",
"sumpmark"
],
"natural/wood":[
"vildmark",
"naturskog",
"skog",
"bush",
"regnskog",
"träd",
"djungel",
"Naturskog",
"urskog"
],
"network/type/node_network":[
"Nod i rekreationsvägsnätverk",
"cykelled",
"vandringsled",
"nodnätverk",
"cykelnätverk",
"vandringsnätverk",
"nod i rekreationsvägsnätverk"
],
"noexit/yes":[
"vägslut",
"återvändsgränd",
"Återvändsgata",
"blindgata återvändsgata"
],
"office":[
"tjänsteman",
"byrå",
"tjänstemän",
"Kontor",
"expedition",
"kontor",
"tjänster"
],
"office/accountant":[
"bokhållare",
"bokföring",
"tjänsteman",
"redovisningsekonom",
"Bokhållare",
"kontorist",
"räkenskap"
],
"office/administrative":[
"Lokal myndighet"
],
"office/adoption_agency":[
"adoption",
"adoptering",
"Adoptionsbyrå",
"barnupptagande",
"adoptionsbyrå",
"adoptera"
],
"office/advertising_agency":[
"Reklambyrå",
"annons",
"annonsbyrå",
"reklam",
"marknadsföring",
"reklambyrå",
"annonsering"
],
"office/architect":[
"arkitektbyrå",
"arkitekt",
"ritningar",
"byggnadskonstnär",
"Arkitektbyrå",
"arkitektkontor",
"byggnadskonst"
],
"office/association":[
"frivillig",
"frivilligorganisation",
"Frivilligorganisation",
"ideell",
"förening",
"volontär",
"organisation",
"frivilligarbetare",
"samhälle",
"icke vinstdrivande",
"biståndsarbetare"
],
"office/bail_bond_agent":[
"bail bond-agent",
"Bail Bond-agent",
"borgen"
],
"office/charity":[
"biståndsorganisation",
"välgörenhet",
"hjälpverksamhet",
"Välgörenhetsorganisation",
"välgörenhetsorganisation",
"bistånd"
],
"office/company":[
"företagskontor",
"expedition",
"kontor",
"Företagskontor",
"kundmottagning",
"företag"
],
"office/consulting":[
"konsultföretag",
"konsulter",
"Konsultkontor",
"konsult",
"konsultkontor"
],
"office/coworking":[
"distansarbete",
"dagkontor",
"kontorsplats",
"coworking",
"mötesrum",
"kontor",
"lånekontor",
"Dagkontor",
"affärslounger",
"tillfällig arbetsplats",
"kontorsarbetsplats",
"tillfälligt kontor",
"fjärrarbetsplats",
"konferensrum"
],
"office/diplomatic":[
"konsulat",
"statssändebud",
"ambassadkontor",
"diplomatkontor",
"diplomat",
"ambassadör",
"envoyé",
"Diplomatkontor",
"ambassad"
],
"office/diplomatic/consulate":[
"konsulat",
"statssändebud",
"ambassadkontor",
"diplomatkontor",
"diplomat",
"ambassadör",
"envoyé",
"ambassad",
"Konsulat"
],
"office/diplomatic/embassy":[
"konsulat",
"statssändebud",
"ambassadkontor",
"diplomatkontor",
"Ambassad",
"diplomat",
"ambassadör",
"envoyé",
"ambassad"
],
"office/diplomatic/liaison":[
"konsulat",
"ambassadkontor",
"diplomatkontor",
"ambassadör",
"envoyé",
"ambassad",
"sambandscentral",
"statssändebud",
"sambandsman",
"kontaktkontor",
"sambandsmän",
"Kontaktkontor",
"diplomat"
],
"office/educational_institution":[
"rektorsexpedition",
"skolledning",
"rektor",
"skolexpedition",
"Utbildningskontor",
"expedition",
"utbildningskontor"
],
"office/employment_agency":[
"förmedling",
"Arbetsförmedling",
"arbetsförmedlingen",
"jobb",
"arbetssökande",
"arbetsförmedling",
"arbetslös"
],
"office/energy_supplier":[
"ström",
"elbolag",
"el",
"gas",
"energibolag",
"Energibolag",
"energi"
],
"office/estate_agent":[
"fastighet",
"husförmedling",
"mäklare",
"fastighetsmäklare",
"fastighetsuthyrning",
"fastighetsförmedling",
"Mäklare/bostadsförmedling",
"egendom",
"bostadsuthyrning",
"bostadsförmedling",
"mark",
"kontorsuthyrning"
],
"office/financial":[
"finans",
"bank",
"bankkontor",
"Bankkontor",
"ekonomisk",
"ekonomi",
"finanskontor"
],
"office/financial_advisor":[
"Finansiell rådgivare",
"arv",
"bankkontor",
"rådgivare",
"sparande",
"kapitalförvaltning",
"ekonomisk",
"finansiell rådgivare",
"aktier",
"finanskontor",
"bank",
"bankman",
"pension",
"ekonomi"
],
"office/forestry":[
"skogsbolag",
"skog",
"skogsvaktare",
"Skogsbolag"
],
"office/foundation":[
"Stiftelse",
"donation",
"stiftelse",
"fond"
],
"office/government":[
"myndighetskontor",
"statlig myndighet",
"Myndighet",
"myndighet"
],
"office/government/prosecutor":[
"åklagarmyndighet",
"åklagare",
"åtal",
"justitieminister",
"Åklagarmyndighet",
"distriktsadvokat"
],
"office/government/register_office":[
"stadshus",
"inskrivningskontor",
"registreringsbyrå",
"folkbokföring",
"registreringskontor",
"mantalslängder",
"skattemyndigheten",
"registrerade enhet",
"Registreringsbyrå",
"borgerlig vigsel"
],
"office/government/tax":[
"Skattekontor",
"skattekontor",
"skattemyndigheten",
"myndighet",
"skatt"
],
"office/guide":[
"rundtur",
"turistguide",
"dykguide",
"Guidekontor",
"guidekontor",
"guide",
"fjällguide"
],
"office/insurance":[
"försäkringar",
"försäkringsförmedling",
"försäkringskontor",
"Försäkringskontor"
],
"office/it":[
"mjukvaruutveckling",
"hårdvara",
"it-specialist",
"IT-kontor",
"it",
"datorer",
"program",
"datorspecialist",
"datakonsult",
"konsultkontor",
"programmering",
"datorkonsult",
"dator",
"it-kontor",
"systemutveckling",
"mjukvara",
"konsult"
],
"office/lawyer":[
"advokat",
"juridiskt ombud",
"jurist",
"lagman",
"rättsombud",
"ombud",
"advokatkontor",
"försvarare",
"Advokatkontor"
],
"office/lawyer/notary":[
"Notariekontor"
],
"office/moving_company":[
"flyttfirma",
"flytt",
"flyttlass",
"Flyttfirma",
"bärare",
"flyttning",
"transport",
"flyttkarl"
],
"office/newspaper":[
"redaktion",
"utgivare",
"nyhetsredaktion",
"tidning",
"Tidningsredaktion",
"tidningslokal",
"magasin",
"tidningsredaktion",
"tidskrift"
],
"office/ngo":[
"frivillig",
"ideell förening",
"icke-statlig organisation",
"frivilligorganisation",
"intresseorganisation",
"ideell",
"förening",
"icke-kommersiell",
"organisation",
"hjälporganisation",
"fackförening",
"Icke-statlig organisation"
],
"office/notary":[
"Notarie",
"arv",
"avtal",
"notarie",
"värdehandlningar",
"bevittna",
"egendom",
"fullmakt",
"handlingar",
"testamente",
"namnteckning",
"notarius",
"notarius publicus",
"dödsbo",
"notariekontor",
"underskrift",
"signatur",
"kontrakt",
"påskrift"
],
"office/physician":[
"Läkare"
],
"office/political_party":[
"Partikontor",
"partihögkvarter",
"partikontor",
"politik",
"parti",
"politiskt parti"
],
"office/private_investigator":[
"detektiv",
"deckare",
"privatdetektiv",
"Privatdetektiv"
],
"office/quango":[
"kvasiautonom",
"Kvasiautonom icke-statlig organisation",
"kvasi",
"organisation",
"quango",
"icke-statlig"
],
"office/religion":[
"religiös",
"församling",
"församlingshem",
"religiöst kontor",
"Religiöst kontor",
"religion"
],
"office/research":[
"efterforskning",
"undersökning",
"forskning",
"utveckling",
"vetenskapligt studium",
"vetenskapligt arbete",
"forskning och utveckling",
"Forskning och utveckling",
"research"
],
"office/security":[
"vakt",
"skyddsvakt",
"säkerhetskontor",
"säkerhetsinspektör",
"Bevakningskontor",
"bevakningskontor",
"väktarkontor",
"områdesbevakning",
"väktare",
"bevakning",
"säkerhetsvakt",
"vaktkontor",
"säkerhet",
"ordningsvakt"
],
"office/surveyor":[
"riskbedömare",
"riskbedömning",
"Undersökning/inspektion",
"inspektion",
"stickprovsundersökning",
"statistik",
"enkät",
"undersökning",
"lantmätare",
"opinionsundersökning",
"skadebedömare",
"skadebedömning",
"lantmäteri",
"mätning"
],
"office/tax_advisor":[
"skatterådgivning",
"ekonomirådgivning",
"skattekonsultation",
"Skatterådgivning",
"skatteplanering",
"moms",
"ekonomi",
"konsultation",
"skatt"
],
"office/telecommunication":[
"mobiltelefon",
"telekom",
"mobiltelefoni",
"surfning",
"internetcafé",
"telefoni",
"telefon",
"Telekom",
"telefoner",
"surfcafé mobil",
"internet"
],
"office/therapist":[
"språkterapi",
"beteendeterapi",
"terapeut",
"fysioterapi",
"kognitiv beteendeterapi",
"psykolog",
"sexterapi",
"kemoterapi",
"samtalsterapi",
"psykologi",
"behandling",
"talterapi",
"cellgiftsbehandling",
"radioterapi",
"röstterapi",
"sjukgymnast",
"farmakoterapi",
"psykoterapi",
"Terapeut",
"familjeterapi",
"behandlare",
"psykoterapeut",
"kognitiv terapi",
"logoped",
"terapi",
"arbetsterapeut",
"psykoanalys",
"arbetsterapi",
"kbt"
],
"office/travel_agent":[
"Resebyrå"
],
"office/water_utility":[
"dricksvatten",
"Vattenleverantör",
"vattenleverantör",
"vattenbolag"
],
"piste/downhill":[
"skidor",
"alpint",
"slalombacke",
"Utförsåkning",
"skidbacke",
"utförsåkning",
"pist",
"snowboard"
],
"piste/downhill/halfpipe":[
"skidor",
"Halfpipe för vintersport",
"alpint",
"skida",
"skidbacke",
"utförsåkning",
"pist",
"vintersport",
"halfpipe",
"half-pipe",
"halfpipe för vintersport",
"slalombacke",
"half pipe",
"snowboard"
],
"piste/hike":[
"vintervandring",
"vandring",
"snöskor",
"skidor",
"Snöskor- / vintervandring",
"vandringsled",
"snöskorvandring",
"pist"
],
"piste/ice_skate":[
"rink",
"skridskorink",
"isbana",
"skridskor",
"skridskoåkning",
"skridskobana",
"Skridskoled",
"is",
"skridskoled",
"pist"
],
"piste/nordic":[
"off-pist",
"längdskidåkning",
"skidor",
"skating",
"skidspår",
"längdåkning",
"pist",
"längdskidor",
"Längdskidspår"
],
"piste/piste":[
"längdskidspår",
"isåkning",
"off-pist",
"vintervandring",
"skridsko",
"alpin",
"skidor",
"utför",
"skidtur",
"släde",
"alpint",
"skida",
"is",
"utförsåkning",
"pist",
"häst",
"längdskidor",
"skidåkning",
"Vintersportspår / Pist",
"vintersportspår",
"snöskor",
"skridskoåkning",
"offpist",
"snowboard"
],
"piste/skitour":[
"skidturåkning",
"skidåkning",
"skidturspår",
"skidtur",
"skidor",
"skidspår",
"Skidturspår",
"pist"
],
"piste/sled":[
"kälke",
"bob",
"rodel",
"släde",
"snowracer",
"pulkabacke",
"pulka",
"Pulkabacke",
"pist"
],
"piste/sleigh":[
"hundspann",
"kälke",
"slädspår",
"husky",
"släde",
"hundsläde",
"Slädspår",
"slädpist",
"pist",
"häst",
"hästsläde"
],
"place":[
"Plats"
],
"place/city":[
"större stad",
"stad",
"metropol",
"storstad",
"världsstad",
"huvudstad",
"Större stad"
],
"place/city_block":[
"bostadskomplex",
"husgrupp",
"kvarter",
"Kvarter"
],
"place/farm":[
"Gård"
],
"place/hamlet":[
"småort",
"gårdar",
"by",
"litet samhälle",
"By",
"gårdssamling"
],
"place/island":[
"holme",
"klippa",
"atoll",
"rev",
"skär",
"ö",
"kobbe",
"Ö",
"skärgård"
],
"place/islet":[
"holme",
"atoll",
"grynna",
"grund",
"rev",
"skär",
"ö",
"kobbe",
"liten ö",
"Holme",
"havsklippa",
"skärgård"
],
"place/isolated_dwelling":[
"bosättning",
"Isolerad boplats",
"isolerad boplats",
"boplats"
],
"place/locality":[
"läge",
"plats",
"lokalitet",
"ställe",
"trakt",
"obefolkad plats",
"Plats"
],
"place/neighbourhood":[
"bostadsområde",
"område",
"närområde",
"kvarter",
"stadsdel",
"Kvarter"
],
"place/plot":[
"lott",
"hustomt",
"tomt",
"privat",
"skifte",
"Tomt",
"trädgård",
"mark"
],
"place/quarter":[
"Kvarter / Under-Borough",
"område",
"kvarter",
"grannskap",
"under-borough",
"stadsdel"
],
"place/square":[
"plaza",
"salutorg",
"marknadsplats",
"torg",
"Torg",
"publik yta",
"stadstorg"
],
"place/suburb":[
"kranskommun",
"förort",
"kommundelsnämnd",
"område",
"stadsområde",
"Förort / Borough",
"förstad",
"kommun",
"grannskap",
"borough",
"stadsdel"
],
"place/town":[
"ort",
"stad",
"Mellanstor stad",
"samhälle"
],
"place/village":[
"ort",
"tätort",
"Mindre samhälle"
],
"playground":[
"Lekplatsutrustning"
],
"playground/balancebeam":[
"Balansbom (lekplats)",
"bom",
"lek",
"lekplats",
"lekområde",
"balansbom",
"balans",
"lekpark"
],
"playground/basketrotator":[
"karusell",
"lek",
"lekplats",
"lekområde",
"korgkarusell",
"lekpark",
"Korgkarusell"
],
"playground/basketswing":[
"lek",
"lekplats",
"lekområde",
"gunga",
"korggunga",
"kompisgunga",
"korg",
"fågelbogunga",
"Korggunga",
"gungställning",
"lekpark"
],
"playground/climbingframe":[
"Klätterställning",
"klättring",
"lek",
"lekplats",
"lekområde",
"klätterställning",
"klättra",
"lekpark"
],
"playground/cushion":[
"Hoppkudde",
"lek",
"lekplats",
"lekområde",
"hoppkudde",
"lekpark"
],
"playground/horizontal_bar":[
"bar",
"lek",
"lekplats",
"lekområde",
"räck",
"lekpark",
"Räck (lekplats)"
],
"playground/playhouse":[
"lek",
"lekplats",
"lekområde",
"Lekhus",
"lekslott",
"lekplatshus",
"lekhus",
"lekstuga",
"lekpark"
],
"playground/roundabout":[
"karusell",
"lek",
"lekplats",
"lekområde",
"Karusell (lekplats)",
"lekpark"
],
"playground/sandpit":[
"sand",
"Sandlåda",
"lek",
"sandlåda",
"lekplats",
"lekområde",
"lekpark"
],
"playground/seesaw":[
"lek",
"gungbräda",
"lekplats",
"lekområde",
"Gungbräda",
"lekpark"
],
"playground/slide":[
"lek",
"lekplats",
"lekområde",
"rutschkana",
"Rutschkana",
"rutschbana",
"lekpark",
"rutchelbana"
],
"playground/springy":[
"lek",
"Fjädergunga",
"lekplats",
"lekområde",
"fjädergunga",
"gungdjur",
"lekpark"
],
"playground/structure":[
"lek",
"lekplats",
"lekområde",
"Lekhus",
"lekslott",
"lekhus",
"lekstuga",
"lekpark"
],
"playground/swing":[
"lek",
"lekplats",
"lekområde",
"gunga",
"Gungställning",
"gungställning",
"lekpark"
],
"playground/zipwire":[
"lek",
"lekplats",
"lekområde",
"Linbana (lekplats)",
"linbana",
"lekpark"
],
"point":[
"läge",
"punkt",
"fläck",
"plats",
"ställe",
"Punkt"
],
"polling_station":[
"val",
"rösta",
"omröstning",
"röstmaskin",
"vallokal",
"valbås",
"valsedel",
"röstning",
"folkomröstning",
"valmaskin",
"Tillfällig vallokal",
"valurna",
"omröstningsapparat"
],
"power":[
"Kraftobjekt"
],
"power/cable":[
"Kraftkabel"
],
"power/cable/underground":[
"kraftledning",
"kraft",
"ström",
"högspänning",
"underjordisk kraftkabel",
"elledning",
"elnät",
"el",
"högspänningsledning",
"strömförsörjning",
"elförsörjning",
"Underjordisk kraftkabel"
],
"power/generator":[
"strömtillverkning",
"Elgenerator",
"kraftgenerator",
"kraftkälla",
"generator",
"elgenerator"
],
"power/generator/method/photovoltaic":[
"solenergi",
"pv-modul",
"fotovoltaik",
"solcell",
"solkraft",
"solljus",
"solkraftverk",
"solpanel",
"termisk solkraft",
"Solpanel",
"solcellsmodul",
"solel"
],
"power/generator/method/photovoltaic/building/roof":[
"soltak",
"solcell",
"solcarport",
"solmarkis",
"solpanel",
"solcellstak",
"Solpaneltak"
],
"power/generator/method/photovoltaic/location/roof":[
"Solpanel på byggnad",
"pv-modul",
"solcell",
"hemsolpanel",
"solpanel",
"taksolcellsmodul",
"taksolpanel"
],
"power/generator/source/hydro":[
"dam",
"vattenkraftverk",
"vattenturbin",
"Vattenkraftverk",
"vattenkraft",
"generator",
"turbin"
],
"power/generator/source/nuclear":[
"kärnanläggning",
"kärnenergi",
"kärnreaktor",
"atomkraftverk",
"kärnkraft",
"kärnkraftsreaktor",
"kärnkraftvärk",
"reaktor",
"atomkraft",
"nukleär energi",
"Kärnkraftsreaktor",
"kärnkraftverk",
"atomenergi",
"kärnkraftsanläggning"
],
"power/generator/source/wind":[
"vindmölla",
"Vindturbin",
"vindturbin",
"vindkraftverk",
"vindkraft"
],
"power/line":[
"kraftledning",
"högspänning",
"elledning",
"högspänningsledning",
"Högspänningsledning"
],
"power/minor_line":[
"kraftledning",
"elledning",
"Mindre kraftledning"
],
"power/plant":[
"el",
"kol",
"generator",
"kraft",
"vind*",
"elkraftverk",
"vattenkraft*",
"kärnkraft*",
"Område för kraftproduktion",
"elproduktion",
"gas",
"solkraft*",
"kraftproduktion"
],
"power/plant/source/coal":[
"kolkraftverk",
"eldkraftverk",
"koleldat kraftverk",
"kraftstation",
"kol",
"fossilkraftverk",
"Koleldat kraftverk",
"fossil"
],
"power/plant/source/gas":[
"gaskraftverk",
"eldkraftverk",
"fossilgas",
"gas",
"kraftstation",
"fossilkraftverk",
"Gaseldat kraftverk",
"fossil",
"gaseldat kraftverk",
"naturgas"
],
"power/plant/source/hydro":[
"dam",
"Vattendrivet kraftverk",
"vattenkraftverk",
"vattenturbin",
"vattenkraft",
"vattendrivet kraftverk",
"vatten",
"turbin"
],
"power/plant/source/nuclear":[
"kärnkraftsverk",
"atomkraft",
"atomkraftverk",
"kraftstation",
"kärnkraft",
"generator",
"Kärnkraftsverk"
],
"power/plant/source/oil":[
"olja",
"eldkraftverk",
"kraftstation",
"fossilkraftverk",
"oljeeldat kraftverk",
"oljekraftverk",
"fossil",
"Oljeeldat kraftverk"
],
"power/plant/source/solar":[
"ljuskraft",
"solpark",
"Solfarm",
"solkraft",
"solkraftverk",
"ljuskraftverk",
"solpanel",
"solfarm"
],
"power/plant/source/waste":[
"avfallsförbränningsanläggning",
"avfall",
"förbränning",
"kraftstation",
"generator",
"sopförbränningsanläggning",
"Avfallsförbränningskraftverk",
"avfallsförbränningskraftverk",
"förgasning",
"avfallsanläggning",
"förbränningsanläggning",
"kraftverk",
"eldkraftverk",
"sopor",
"graftverk"
],
"power/plant/source/wind":[
"vindfarm",
"vindpark",
"vindmölla",
"Vindfarm",
"vindturbin",
"vindkraftverk",
"vindkraft",
"vind"
],
"power/pole":[
"elledningsstolpe",
"mast",
"stolpe",
"Kraftledningsstolpe",
"kraftledningsstolpe",
"kraftledningsmast",
"elledningsmast"
],
"power/substation":[
"elomvandling",
"transformator",
"Fördelningsstation",
"fördelningsstation",
"stadsnätstation",
"elskåp",
"elfördelning"
],
"power/switch":[
"frånskiljare",
"Frånskiljare",
"strömbrytare"
],
"power/tower":[
"mast",
"högspänningsmast",
"Högspänningsmast",
"kraftledningsstolpe",
"kraftledningsmast"
],
"power/transformer":[
"elomvandling",
"transformator",
"nätstation",
"Transformator"
],
"public_transport/platform":[
"väntplats",
"kollektivtrafik",
"transit",
"avsats",
"plattform",
"Plattform för kollektivtrafik",
"transport",
"påstigningsplats",
"perrong"
],
"public_transport/platform/aerialway":[
"Linbaneplattform",
"linbanestopp",
"hållplats",
"stopp",
"linbaneterminal",
"aerialway",
"linbana",
"terminal",
"linjetrafik",
"transport",
"linbanehållplats",
"kollektivtrafik",
"transit",
"plattform",
"linbaneplattform"
],
"public_transport/platform/aerialway_point":[
"Hållplats / Plattform för linbana"
],
"public_transport/platform/bus":[
"busshållplats",
"kollektivtrafik",
"hållplats",
"bussplattform",
"Bussplattform",
"transit",
"plattform",
"transport",
"linjetrafik",
"buss"
],
"public_transport/platform/bus_point":[
"Busshållplats",
"busshållplats",
"busstation",
"hållplats",
"station",
"busstopp",
"anhalt",
"buss"
],
"public_transport/platform/bus_tram_point":[
"busshållplats",
"busstation",
"hållplats",
"spårvägshållplats",
"spårvagnstopp",
"anhalt",
"spårvagns- & busstopp",
"Spårvagns- & busstopp",
"spårväg",
"kollektivtrafik",
"spårvagnsterminal",
"spårvagn",
"station",
"plattform",
"spårvagnshållplats",
"busstopp",
"spår",
"buss"
],
"public_transport/platform/ferry":[
"färjestation",
"brygga",
"färjehållplats",
"stopp",
"färjeterminal",
"båthållplats",
"färjestopp",
"terminal",
"linjetrafik",
"transport",
"färja",
"båt",
"färjeplattform",
"kollektivtrafik",
"båtterminal",
"Färjeplattform",
"transit",
"pir",
"station",
"plattform",
"båtstopp"
],
"public_transport/platform/ferry_point":[
"Stop / plattform för färja"
],
"public_transport/platform/light_rail":[
"Hållplats för snabbspårväg / stadsbana",
"hållplats",
"light rail",
"spårvagnsplattform",
"vagn",
"spårvägshållplats",
"stadsbana",
"terminal",
"transport",
"snabbspårväg",
"spårväg",
"kollektivtrafik",
"spårvagnsterminal",
"transit",
"spårvagn",
"plattform",
"järnväg",
"spår"
],
"public_transport/platform/light_rail_point":[
"Hållplats för snabbspårväg / stadsbana"
],
"public_transport/platform/monorail":[
"monorailstopp",
"stopp",
"Plattform för monorail",
"enskensbana",
"linjetrafik",
"transport",
"räls",
"monorail",
"monorailplattform",
"kollektivtrafik",
"plattform",
"balkbana",
"spår"
],
"public_transport/platform/monorail_point":[
"Stopp / plattform för monorail"
],
"public_transport/platform/subway":[
"Tunnelbaneplattform",
"kollektivtrafik",
"metro",
"tunnelbanestopp",
"plattform",
"transport",
"tunnelbana",
"järnväg",
"spår",
"underjordisk",
"tunnelbaneplattform"
],
"public_transport/platform/subway_point":[
"Tunnelbanestopp / -plattform"
],
"public_transport/platform/train":[
"järnvägsperrong",
"stopp",
"järnvägsplattform",
"linjetrafik",
"transport",
"tågstopp",
"kollektivtrafik",
"transit",
"tåg",
"Järnvägsperrong",
"plattform",
"perrong",
"järnväg",
"spår"
],
"public_transport/platform/train_point":[
"Järnvägsstopp / -perrong"
],
"public_transport/platform/tram":[
"hållplats",
"spårvagnsplattform",
"vagn",
"spårvägshållplats",
"Spårvagnsplattform",
"terminal",
"transport",
"spårväg",
"kollektivtrafik",
"spårvagnsterminal",
"transit",
"spårvagn",
"plattform",
"spårvagnshållplats",
"järnväg"
],
"public_transport/platform/tram_point":[
"hållplats",
"spårvagnsplattform",
"vagn",
"spårvägshållplats",
"Spårvagnshållplats / -plattform",
"terminal",
"transport",
"spårväg",
"kollektivtrafik",
"spårvagnsterminal",
"transit",
"spårvagn",
"plattform",
"spårvagnshållplats",
"järnväg"
],
"public_transport/platform/trolleybus":[
"busshållplats",
"hållplats",
"spårlös",
"vagn",
"transport",
"trådbuss",
"kollektivtrafik",
"bussplattform",
"transit",
"spårvagn",
"plattform",
"Bussplattform för trådbuss",
"buss"
],
"public_transport/platform/trolleybus_point":[
"busshållplats",
"hållplats",
"spårlös",
"vagn",
"transport",
"trådbuss",
"kollektivtrafik",
"bussplattform",
"transit",
"spårvagn",
"plattform",
"Busshållplats för trådbuss",
"buss"
],
"public_transport/platform_point":[
"väntplats",
"avsats",
"plattform",
"Hållplats / Plattform för kollektivtrafik",
"påstigningsplats",
"perrong"
],
"public_transport/station":[
"kollektivtrafik",
"Station för kollektivtrafik",
"bytespunkt",
"station",
"resecenter",
"station för kollektivtrafik",
"terminal",
"transport"
],
"public_transport/station_aerialway":[
"linbanestation",
"kollektivtrafik",
"transit",
"station",
"aerialway",
"Linbanestation",
"linbana",
"terminal",
"transport"
],
"public_transport/station_bus":[
"busshållplats",
"busstation",
"kollektivtrafik",
"bussterminal",
"transit",
"station",
"resecenter",
"reseterminal",
"terminal",
"transport",
"Busstation / Bussterminal",
"buss"
],
"public_transport/station_ferry":[
"färjestation",
"brygga",
"färjehållplats",
"färjeterminal",
"båthållplats",
"Färjeterminal",
"terminal",
"transport",
"färja",
"båt",
"kollektivtrafik",
"båtterminal",
"transit",
"pir",
"station"
],
"public_transport/station_light_rail":[
"light rail",
"lättbana",
"hållplats",
"station för snabbspårväg",
"stadsbana",
"spårvagnstopp",
"Station för snabbspårväg / stadsbana",
"transport",
"linjetrafik",
"terminal",
"snabbspårväg",
"spårväg",
"kollektivtrafik",
"spårvagnsterminal",
"station för light rail",
"spårvagn",
"station",
"spårvagnshållplats",
"järnväg",
"spår"
],
"public_transport/station_monorail":[
"enskensbana",
"terminal",
"linjetrafik",
"transport",
"monorailstation",
"räls",
"monorail",
"kollektivtrafik",
"station",
"plattform",
"Monorailstation",
"spår",
"balkbana"
],
"public_transport/station_subway":[
"tunnelbanestation",
"kollektivtrafik",
"metro",
"station",
"transport",
"terminal",
"tunnelbana",
"järnväg",
"spår",
"underjordisk",
"Tunnelbanestation"
],
"public_transport/station_train":[
"linjeplats",
"trafikplats",
"central",
"tåghållplats",
"hållplats",
"järnvägshållplats",
"Järnvägsstation",
"centralstation",
"huvudbangård",
"hållställe",
"järnvägsstation",
"tågstation"
],
"public_transport/station_train_halt":[
"hållplats",
"hållställe",
"transport",
"avstigning",
"Mindre järnvägshållplats",
"kollektivtrafik",
"järnvägshållplats",
"påstigning",
"transit",
"tåg",
"station",
"plattform",
"järnvägsstation",
"järnväg",
"spår",
"mindre järnvägshållplats"
],
"public_transport/station_tram":[
"spårväg",
"Spårvagnsstation",
"spårvagnsterminal",
"spårvagn",
"station",
"spårvägshållplats",
"spårvagnsstation"
],
"public_transport/station_trolleybus":[
"busshållplats",
"hållplats",
"station / terminal för trådbuss",
"terminal",
"linjetrafik",
"transport",
"Station / Terminal för trådbuss",
"trådbussterminal",
"trådbuss",
"trådbusstopp",
"kollektivtrafik",
"bussterminal",
"station",
"busstopp",
"trådbusshållplats",
"buss"
],
"public_transport/stop_area":[
"kollektivtrafik",
"hållplats",
"bytespunkt",
"transit",
"byte",
"station",
"knutpunkt",
"resecenter",
"terminal",
"linjetrafik",
"transport",
"Bytespunkt / knutpunkt"
],
"public_transport/stop_position":[
"stopposition för kollektivtrafik",
"stopposition",
"kollektivtrafik",
"hållplats",
"Stopposition för kollektivtrafik",
"linjetrafik",
"transport"
],
"public_transport/stop_position_aerialway":[
"stopposition",
"Stopposition för linbana",
"linbanestation",
"linbanestopp",
"stopposition för linbana",
"kollektivtrafik",
"hållplats",
"linbaneterminal",
"linbana",
"linjetrafik",
"transport",
"linbanehållplats"
],
"public_transport/stop_position_bus":[
"stopposition för buss",
"stopposition",
"busshållplats",
"kollektivtrafik",
"hållplats",
"bussterminal",
"busstopp",
"linjetrafik",
"transport",
"buss",
"Stopposition för buss"
],
"public_transport/stop_position_ferry":[
"båt",
"stopposition",
"busshållplats",
"stopposition för färja",
"kollektivtrafik",
"hållplats",
"bussterminal",
"busstopp",
"linjetrafik",
"transport",
"färja",
"Stopposition för färja"
],
"public_transport/stop_position_light_rail":[
"stopposition",
"light rail",
"lättbana",
"hållplats",
"stadsbana",
"spårvagnstopp",
"transport",
"linjetrafik",
"snabbspårväg",
"spårväg",
"kollektivtrafik",
"spårvagnsterminal",
"spårvagn",
"Stopposition för snabbspårväg / stadsbana",
"spårvagnshållplats",
"järnväg",
"spår",
"stopposition för snabbspårväg"
],
"public_transport/stop_position_monorail":[
"stopposition",
"kollektivtrafik",
"hållplats",
"Stopposition för monorail",
"enskensbana",
"linjetrafik",
"transport",
"balkbana",
"spår",
"stopposition för monorail",
"räls",
"monorail"
],
"public_transport/stop_position_subway":[
"tunnelbanetåg",
"stopposition",
"tunnelbanestation",
"kollektivtrafik",
"hållplats",
"tunnelbanestopp",
"stopposition för tunnelbana",
"linjetrafik",
"transport",
"tunnelbana",
"tunnelbanehållplats",
"Stopposition för tunnelbana"
],
"public_transport/stop_position_train":[
"tågterminal",
"järnvägsstopp",
"stopposition",
"hållplats",
"linjetrafik",
"transport",
"tågstopp",
"kollektivtrafik",
"järnvägshållplats",
"tåg",
"järnvägsterminal",
"stopposition för tåg",
"järnvägsstation",
"tågstation",
"Stopposition för tåg"
],
"public_transport/stop_position_tram":[
"stopposition",
"kollektivtrafik",
"hållplats",
"spårvagnsterminal",
"spårvagn",
"Stopposition för spårvagn",
"spårvagnstopp",
"spårvagnshållplats",
"linjetrafik",
"transport",
"stopposition för spårvagn"
],
"public_transport/stop_position_trolleybus":[
"stopposition",
"busshållplats",
"hållplats",
"Stopposition för trådbuss",
"linjetrafik",
"transport",
"trådbussterminal",
"stopposition för trådbuss",
"trådbuss",
"trådbusstopp",
"kollektivtrafik",
"bussterminal",
"busstopp",
"trådbusshållplats",
"buss"
],
"railway":[
"Järnvägsobjekt"
],
"railway/abandoned":[
"borttagen järnväg",
"riven järnväg",
"Uppriven spårsträcka"
],
"railway/buffer_stop":[
"Stoppbock",
"stoppbock",
"buffert",
"buffertstopp",
"stoppblock"
],
"railway/construction":[
"järnväg under uppförande",
"bygge",
"Spår under uppbyggnad",
"byggarbete",
"byggnadsplats",
"järnväg under byggnad",
"järnväg under konstruktion",
"järnväg",
"byggarbetsplats",
"byggnation"
],
"railway/crossing":[
"spårpassage",
"järnvägspassage",
"cykelväg",
"gångväg",
"stig",
"tågkorsning",
"plankorsning",
"tågövergång",
"cykelpassage",
"Järnvägskorsning (stig)",
"gångpassage",
"järnvägskorsning",
"tågpassage",
"korsning",
"järnvägsövergång",
"övergångsställe"
],
"railway/derail":[
"utspårare",
"Spårspärr",
"omläggningsanordning",
"spårspärr"
],
"railway/disused":[
"övergiven järnväg",
"Nedlagd spårsträcka",
"oanvänd tågbana",
"oanvänd järnväg",
"övergiven tågbana"
],
"railway/funicular":[
"bergbana",
"klippbana",
"linbana",
"Bergbana"
],
"railway/halt":[
"Mindre järnvägshållplats"
],
"railway/level_crossing":[
"spårpassage",
"järnvägspassage",
"tågkorsning",
"plankorsning",
"tågövergång",
"järnvägskorsning",
"Järnvägskorsning (väg)",
"tågpassage",
"korsning",
"järnvägsövergång"
],
"railway/light_rail":[
"smalspår",
"smalspårig järnväg",
"Snabbspårväg / stadsbana",
"stadsbana",
"järnväg",
"snabbspårväg"
],
"railway/milestone":[
"kilometertavla",
"kilometerpåle",
"milsten",
"referenstavla",
"kilometerstolpe",
"Kilometerstolpe vid järnväg",
"avståndsmärke"
],
"railway/miniature":[
"smalspår",
"smalspårig järnväg",
"trädgårdsjärnväg",
"miniatyrjärnväg",
"Miniatyrjärnväg",
"åkbar miniatyrjärnväg"
],
"railway/monorail":[
"Monorail",
"kollektivtrafik",
"enskensbana",
"linjetrafik",
"transport",
"balkbana",
"spår",
"räls",
"monorail"
],
"railway/monorail/hanging":[
"hängande enskensbana",
"hängande monorail-spår",
"hängande balkbana",
"hängande järnväg",
"Hängande monorail-spår"
],
"railway/narrow_gauge":[
"smalspårig bana",
"smalspår",
"smalspårig järnväg",
"Smalspårbana",
"smalspårig",
"smalspårbana",
"järnväg"
],
"railway/platform":[
"Järnvägsperrong"
],
"railway/preserved":[
"historisk järnväg",
"museijärnväg",
"historiskt tåg",
"turistjärnväg",
"turisttåg",
"Museijärnväg",
"bevarad järnväg",
"ångtåg"
],
"railway/rail":[
"järnvägsspår",
"Järnväg",
"spår",
"bana",
"räls"
],
"railway/rail/highspeed":[
"höghastighetsbana",
"snabbspår",
"järnvägsspår",
"snabbjärnväg",
"höghastighet",
"järnväg",
"spår",
"bana",
"Höghastighetsbana",
"räls"
],
"railway/railway_crossing":[
"spårkors",
"tågkorsning",
"plankorsning",
"korsande järnvägsspår",
"järnvägskorsning",
"korsning",
"Korsning järnväg/järnväg",
"järnväg-järnvägskorsning",
"spårkryss",
"diamantkorsning"
],
"railway/signal":[
"semafor",
"huvudsignal",
"järnvägssignal",
"järnvägsljus",
"försignal",
"signal",
"ljus",
"Järnvägssignal",
"dvärgsignal"
],
"railway/station":[
"Järnvägsstation"
],
"railway/subway":[
"t-bana",
"tunnelbanespår",
"metro",
"underjordisk järnväg",
"tunnelbana",
"Tunnelbana"
],
"railway/subway_entrance":[
"tunnelbaneingång",
"Tunnelbaneingång",
"t-banenedgång",
"t-baneingång",
"tunnelbanenergång"
],
"railway/switch":[
"korsningsväxel",
"järnvägskorsning",
"växel",
"Järnvägsväxel",
"korsning",
"järnvägsväxel"
],
"railway/train_wash":[
"tvätthall",
"tågtvätt",
"Tågtvätt",
"loktvätt"
],
"railway/tram":[
"spårvägsspår",
"spårväg",
"motorvagn",
"spårvagn",
"Spårväg"
],
"railway/tram_crossing":[
"spårvagnskorsning",
"korsande spårvagnsspår",
"plankorsning",
"korsande spårvägsspår",
"korsning",
"korsande",
"spårvägsskorsning",
"Korsning spårvagn/gångväg"
],
"railway/tram_level_crossing":[
"spårvagnskorsning",
"korsande spårvagnsspår",
"plankorsning",
"korsande spårvägsspår",
"korsning",
"Korsning spårvagn/väg",
"korsande",
"spårvägsskorsning"
],
"railway/tram_stop":[
"Stopposition för spårvagn"
],
"railway/yard":[
"rangerbangård",
"godsvagnstopp",
"godstågstation",
"bangård",
"växlingsbangårdar",
"järnvägsstation",
"järnvägsgård",
"kombiterminal",
"Bangård",
"godsbangård"
],
"relation":[
"Relation",
"samband",
"relaterat",
"koppling",
"anknytning",
"förbindelse",
"förhållande",
"kontext",
"relation"
],
"route/ferry":[
"färjelinje",
"båtlinje",
"båtrutt",
"rutt",
"färja",
"Färjerutt",
"färjerutt",
"båt i linjetrafik"
],
"seamark":[
"Sjömärke"
],
"seamark/beacon_isolated_danger":[
"Punktmärke",
"punktmärke",
"iala"
],
"seamark/beacon_lateral":[
"fastmärke",
"farledsmärke",
"lateralmärke",
"iala",
"Farledsmärke",
"farled"
],
"seamark/buoy_lateral":[
"Farledsboj",
"farledsboj",
"farledsmärke",
"lateralmärke",
"boj",
"farled",
"lateralboj"
],
"seamark/buoy_lateral/green":[
"Grön prick",
"grön boj",
"lateralmärke",
"flytande styrbordsmärke",
"iala",
"grön prick",
"styrbordsmärke"
],
"seamark/buoy_lateral/red":[
"röd boj",
"lateralmärke",
"Röd prick",
"röd prick",
"flytande babordsmärke",
"babordsmärke"
],
"seamark/mooring":[
"knap",
"krysshult",
"förtöjningspåle",
"påle",
"förtöjning",
"Förtöjning",
"boj",
"pollare"
],
"shop":[
"shop",
"butik",
"affär",
"Affär"
],
"shop/agrarian":[
"jordbruksmaskiner",
"Jordbruksaffär",
"djurmat",
"jordbruksaffär",
"utsäde",
"frön",
"jordbruk",
"gödsel",
"gödningsmedel",
"jordbruksverktyg",
"lantmannaföreningen",
"bekämpningsmedel",
"jordbruksutrustning"
],
"shop/alcohol":[
"vinaffär",
"spritaffär",
"systemet",
"öl",
"systembolaget",
"Vin-och-spritaffär",
"bolaget",
"vin- och spritaffär",
"alkohol",
"sprit",
"vin- och sprit",
"vin"
],
"shop/anime":[
"cosplay",
"anime/manga-affär",
"figurer",
"japan",
"manga",
"dakimakura",
"Anime/Manga-affär",
"anime"
],
"shop/antiques":[
"antikvitetsaffär",
"antikt",
"antikshop",
"Antikaffär",
"antikvariat",
"antikaffär"
],
"shop/appliance":[
"tvättmaskin",
"vitvarukedja",
"vitvaruaffär",
"mikrovågsugn",
"köksfläkt",
"spis",
"frys",
"hushållsmaskin",
"Vitvaror",
"hushållsmaskiner",
"kylskåp",
"ugn",
"vitvaror",
"vitvara",
"diskmaskin"
],
"shop/art":[
"konstaffär",
"konstverk",
"Konstaffär",
"tavlor",
"kulturer",
"konst",
"konsthandlare",
"konstgalleri",
"galleri",
"statyer",
"konstutställning"
],
"shop/baby_goods":[
"nappflaskor",
"bäbis",
"nappar",
"babykläder",
"spjälsängar",
"Babyprodukter",
"småbarn",
"babyprodukter",
"baby",
"barnkläder",
"bäbiskläder",
"barnvagnar",
"blöjor"
],
"shop/bag":[
"bagageväskor",
"resväskor",
"bagage",
"handväska",
"väskor",
"väskaffär",
"plånbok",
"Väskaffär",
"handväskor"
],
"shop/bakery":[
"bröd",
"Bageri",
"bageri",
"bullar",
"baka",
"bagare"
],
"shop/bathroom_furnishing":[
"Badrumsinredning",
"badrum",
"badrumsinredning"
],
"shop/beauty":[
"Skönhetssalong",
"nagelsalong",
"spa",
"skönhetssalong",
"skönhet",
"kuranstalt",
"smink",
"salong",
"kosmetik",
"solarium",
"shiatsu",
"hälsoanläggning",
"kurort",
"naglar",
"skönhetsbehandlingar",
"massage"
],
"shop/beauty/nails":[
"nagel",
"nagelvård",
"nagelsalong",
"naglar",
"manikur",
"handvård",
"händer",
"manikyr",
"Nagelsalong",
"pedikyr",
"hand",
"manikyrist  manikyrera"
],
"shop/beauty/tanning":[
"solarium",
"konstgjort solljus",
"Solarium"
],
"shop/bed":[
"sängaffär",
"madrasser",
"sängar",
"påslakan",
"Sängaffär",
"täcken",
"lakan",
"kuddar"
],
"shop/beverages":[
"dricka",
"läsk",
"dryck",
"alkohol",
"Dryckaffär",
"läskedryck"
],
"shop/bicycle":[
"cykelförsäljning",
"Cykelaffär",
"cykelaffär",
"cykel",
"cykelreparatör"
],
"shop/boat":[
"båttillbehör",
"båtaffär",
"motorboat",
"Båtaffär",
"båt",
"fiskebåt",
"vattenskoter",
"roddbåt",
"segelbåt",
"segel",
"eka",
"jet-ski",
"jetski"
],
"shop/bookmaker":[
"spel",
"måltipset",
"trav",
"vadslagning",
"dobbel",
"Vadslagning",
"vadhållning",
"stryktipset"
],
"shop/books":[
"Bokhandel",
"bokhandel",
"antikvariat",
"bokförsäljning"
],
"shop/boutique":[
"Boutique (Dyra kläder och accessoarer)"
],
"shop/brewing_supplies":[
"bryggning",
"vintillverkning",
"Affär för hembryggningstillbehör",
"öl",
"vinbryggning",
"affär för hembryggningstillbehör",
"hembryggning",
"vin",
"öltillverkning",
"ölbryggning"
],
"shop/butcher":[
"Slaktare",
"köttaffär",
"charkuterihandlare",
"chark",
"köttstyckare",
"slaktare",
"styckare",
"kött",
"charkuterist"
],
"shop/camera":[
"fotografering",
"Affär för kameratillbehör",
"foto",
"kameratillbehör. kamera",
"linser",
"kameratillbehöraffär",
"film",
"objektiv",
"affär för kameratillbehör"
],
"shop/candles":[
"värmeljus",
"Ljusaffär",
"ljusaffär",
"mysljus",
"ljusstakar",
"ljus",
"stearinljus"
],
"shop/cannabis":[
"420",
"cannabisaffär",
"pot",
"reefer",
"Cannabisaffär",
"cannabis",
"marijuana",
"weed"
],
"shop/car":[
"bilfirma",
"bilhandlare",
"bilreparatör",
"bilförsäljning",
"bilverkstad",
"bilsäljare",
"biltillbehör",
"Bilhandlare"
],
"shop/car/second_hand":[
"bilar",
"bilhandlare med begagnade bilar",
"begagnat",
"begagnade bilar",
"Bilhandlare med begagnade bilar"
],
"shop/car_parts":[
"bilreservdelar",
"motor",
"Biltillbehör",
"bildelar",
"reservdelar",
"biltillbehör"
],
"shop/car_repair":[
"motor",
"bilreparatör",
"Bilverkstad",
"bilverkstad",
"verkstad"
],
"shop/caravan":[
"tältvagn",
"husvagnsförsäljare",
"husbil",
"husvagn",
"husbilsförsäljare",
"Husvagnsförsäljare"
],
"shop/carpet":[
"matta",
"Mattaffär",
"mattaffär",
"mattor"
],
"shop/catalogue":[
"katalog",
"katalogaffär",
"Katalogaffär"
],
"shop/charity":[
"myrorna",
"begagnat",
"secondhandbutik",
"välgörenhetsbutik",
"andrahandsbutik",
"second hand",
"secondhand",
"second hand-butik",
"begagnade varor",
"bättre begagnat",
"vintage",
"Second hand-butik",
"second handbutik",
"välgörenhet"
],
"shop/cheese":[
"ost",
"ostar",
"ostaffär",
"Ostaffär",
"ostbutik"
],
"shop/chemist":[
"hygienartiklar",
"kosmetik",
"kemi",
"kemiaffär",
"städ",
"rengöring",
"smink",
"hygien",
"kosmetika",
"städmaterial",
"Kemiaffär (hygien,  kosmetika & städ)",
"rengöringsmedel"
],
"shop/chocolate":[
"pralin",
"konfekt",
"choklad",
"Chokladaffär",
"chokladaffär",
"praliner"
],
"shop/clothes":[
"klädbutik",
"ekipering",
"Klädaffär",
"klädaffär",
"kläder"
],
"shop/clothes/second_hand":[
"klädbutik",
"klänningar",
"secondhandkläder",
"kostymer",
"Affär med secondhandkläder",
"kjolar",
"begagnade",
"secondhand",
"affär för secondhandkläder",
"skjortor",
"byxor",
"blusar",
"shorts",
"kläder"
],
"shop/clothes/underwear":[
"mode",
"Underklädersaffär",
"kalsonger",
"bh",
"underklänning",
"underkläder",
"trosor",
"lingeri",
"strumpor",
"damunderkläder",
"underklädersaffär",
"sockar"
],
"shop/clothes/wedding":[
"festkläder",
"affär med bröllopskläder",
"brud",
"Affär med bröllopskläder",
"brudtärna",
"bröllopsklänning",
"smoking",
"brudklänning",
"brudgum",
"frack",
"bröllop"
],
"shop/coffee":[
"kaffeaffär",
"kaffepulver",
"Kaffeaffär",
"kaffeböner",
"kaffebönor",
"bryggkaffe",
"kaffe"
],
"shop/collector":[
"mynt",
"samlare",
"medaljer",
"figurer",
"Affär med samlarobjekt",
"samling",
"affär med samlarobjekt",
"serier",
"filateli",
"dockor",
"frimärken'",
"numismatik",
"antikviteter"
],
"shop/computer":[
"data",
"dator",
"datorbutik",
"datorförsäljning",
"Datorbutik",
"datorer",
"datoraffär",
"datorhårdvara",
"datorprogram"
],
"shop/confectionery":[
"konfektyr",
"choklad",
"sötsaker",
"godisbutik",
"godisaffär",
"godis",
"Godisaffär",
"konfektbutik",
"karameller"
],
"shop/convenience":[
"närbutik",
"livsmedelsbutik",
"mataffär",
"Närbutik",
"kvartersbutik",
"livsmedel"
],
"shop/copyshop":[
"kopiering",
"Tryckeri",
"tryckeri",
"copyshop"
],
"shop/cosmetics":[
"sminkaffär",
"Sminkaffär",
"smink",
"kosmetika",
"kosmetikaffär"
],
"shop/country_store":[
"lanthandel",
"Lanthandel",
"landet"
],
"shop/craft":[
"konstverk",
"hantverk",
"konsthantverk",
"konst",
"Konst- & hantverksbutik",
"slöjd"
],
"shop/curtain":[
"Gardinaffär",
"drapera",
"fönster",
"draperier",
"gardiner",
"gardinaffär"
],
"shop/dairy":[
"ost",
"mejeriaffär",
"ägg",
"mejeri",
"mjölk",
"mjölkaffär",
"Mejeriaffär"
],
"shop/deli":[
"lunch",
"smörgås",
"delikatessaffär",
"delikatess",
"Delikatessaffär",
"delikatesser",
"finmat",
"kött"
],
"shop/department_store":[
"Varuhus",
"varuhus",
"affärshus"
],
"shop/doityourself":[
"indie",
"handverktyg",
"heminredning",
"elverktyg",
"byggvaruhus",
"byggmarknad",
"inredning",
"byggsatser",
"verktyg",
"byggsats",
"gördetsjälv",
"gör-det-själv",
"gör det själv",
"Byggmarknad",
"byggmaterial",
"järnaffär",
"bygghandel"
],
"shop/doors":[
"affär med dörrar",
"dörr",
"dörreparation",
"Affär med dörrar",
"dörrar",
"dörrepatör",
"dörrförsäljning"
],
"shop/dry_cleaning":[
"kemtvättar",
"Kemtvätt",
"kemisk tvätt"
],
"shop/e-cigarette":[
"elektrisk cigarett",
"elcigarett",
"Affär för elektroniska cigaretter",
"e-cigarett",
"affär för elektroniska cigaretter"
],
"shop/electrical":[
"kabel",
"el",
"kablage",
"elutrustning",
"kablar",
"led",
"amatur",
"kraft",
"affär med elutrustning",
"fläkt",
"Affär med elutrustning",
"elektronik",
"belysning"
],
"shop/electronics":[
"elektronikbutik",
"spisar",
"tv",
"batterier",
"tvättmaskin",
"kablar",
"datorer",
"radio",
"apparater",
"dator",
"hemelektronik",
"kylskåp",
"torktumlare",
"vitvaror",
"Elektronikbutik",
"hushållsapparater",
"ljud"
],
"shop/erotic":[
"erotik",
"sexaffär",
"sex",
"sexleksaker",
"sexshop",
"porr",
"pornografi",
"porrfilmer",
"Sexshop",
"erotikaffär",
"porrtidningar",
"underkläder",
"sexfilmer",
"kondomer",
"erotisk"
],
"shop/erotic/lgbtq":[
"erotik",
"sexaffär",
"lesbisk",
"sex",
"hbtq",
"sexleksaker",
"sexshop",
"porr",
"pornografi",
"porrfilmer",
"erotikaffär",
"porrtidningar",
"underkläder",
"hbtq-sexshop",
"sexfilmer",
"kondomer",
"gay",
"HBTQ-sexshop",
"erotisk"
],
"shop/fabric":[
"tyg",
"Tygaffär",
"tyger",
"sy",
"tygaffär",
"sömnad"
],
"shop/farm":[
"närproducerat",
"gårdsbutik",
"Gårdsbutik",
"egenproducerat"
],
"shop/fashion":[
"Modebutik"
],
"shop/fashion_accessories":[
"plånböcker",
"Affär för modeaccessoarer",
"affär för modeaccessoarer",
"paraply",
"klockor",
"handväskor",
"modeaccessoarer",
"solglasögon",
"hattar",
"parfym",
"smycken",
"doft",
"väskor",
"accessoarer",
"halsdukar"
],
"shop/fireplace":[
"kakelugn",
"eldstad",
"Kaminbutik",
"gaskamin",
"eldstäder",
"kamin"
],
"shop/fishing":[
"fiskeutrustning",
"vinterfiske",
"fiskeaffär",
"fiske",
"fisk",
"sommarfiske",
"levande bete",
"fiskare",
"fiska",
"bete",
"Fiskeaffär"
],
"shop/flooring":[
"golv",
"parkett",
"klinkergolv",
"golvläggning",
"Affär för golv"
],
"shop/florist":[
"bukett",
"Florist",
"blomsterhandlare",
"blommor",
"florist",
"blomsterbindare",
"blomförsäljning"
],
"shop/frame":[
"Ramaffär",
"ramaffär",
"ramar",
"inramning"
],
"shop/frozen_food":[
"färdigmat",
"mat",
"fryst mat",
"färdigrätter",
"lunch",
"matlådor",
"frys",
"snabbmat",
"frysmat",
"färdigrätt",
"Affär för fryst mat",
"fryst"
],
"shop/fuel":[
"fotogen",
"Bränsleaffär",
"lpg",
"träkol",
"bränslebutik",
"eldningsolja",
"bränsle",
"kol",
"propan",
"bränsleaffär",
"motorbränsle"
],
"shop/funeral_directors":[
"gravsten",
"bodelning",
"begravning",
"jordfästning",
"gravsättning",
"begravningsentreprenör",
"Begravningsbyrå",
"kremering",
"begravningsbyrå",
"gravstenar",
"begravningsceremoni"
],
"shop/furniture":[
"möbelgrossist",
"bord",
"hylla",
"soffor",
"inredning",
"stol",
"stolar",
"Möbelaffär",
"möbelaffär",
"möbelvaruhus",
"soffa"
],
"shop/games":[
"affär för brädspel",
"tärningsspel",
"spelbutik",
"spel",
"live action-rollspel",
"brädspel",
"Affär för brädspel",
"kortspel",
"strategispel",
"miniatyrer krigsspel"
],
"shop/garden_centre":[
"krukväxter",
"trädgårdsväxter",
"jord",
"Trädgårdscenter",
"träd",
"trädgårdsverktyg",
"trädgårdscenter",
"planteringsjord",
"kompost",
"blomkrukor",
"blommor",
"landskap",
"plantskola",
"buskar",
"trädgård"
],
"shop/gas":[
"gasbehållare",
"lpg",
"metangas",
"gasflaskor",
"propan",
"Försäljning av gas",
"naturgas",
"gasol",
"fordonsgas",
"återfyllning",
"gas",
"cng",
"gasolflaskor"
],
"shop/general":[
"generell affär",
"byaffär",
"Generell affär"
],
"shop/gift":[
"presentbutik",
"gratulationskort",
"souvenirbutik",
"grattiskort",
"presenter",
"souvenirer",
"gåva",
"present",
"Presentbutik",
"gåvor",
"souvenir"
],
"shop/greengrocer":[
"frukt",
"frukthandlare",
"grönsaker",
"frukthandel",
"grönsakshandlare",
"Grönsakshandlare",
"vegetabiliskt"
],
"shop/hairdresser":[
"hårfrisör",
"hårkonstnär",
"skägg",
"skönhet",
"skönhetssalong",
"hårförlängning",
"hårkreatör",
"salong",
"stylist",
"hårklippning",
"barberare",
"rakning",
"frisör",
"hår",
"hårtvätt",
"hårfärgning",
"Hårfrisör"
],
"shop/hairdresser_supply":[
"schampo",
"frisör",
"hårspray",
"balsam",
"skönhetsmedel",
"konstgjorda naglar",
"frisyr",
"frisörtillbehör",
"hårförlängningar",
"Affär för hårprodukter"
],
"shop/hardware":[
"handverktyg",
"nycklar",
"spik",
"järntillbehör",
"hushållsprodukter",
"redskap",
"Järnaffär",
"metallverktyg",
"bultar",
"bygg",
"lås",
"järnaffär",
"kök",
"elverktyg",
"badrum",
"krokar",
"el",
"verktyg",
"skruvar",
"trädgårdsredskap",
"nyckeltillverkning",
"vvs",
"järnhandlare",
"bult",
"järnbeslag",
"köksutrustning",
"skruv"
],
"shop/health_food":[
"Hälsokostbutik",
"kosttillskott",
"naturligt",
"organisk",
"vegan",
"mjölkersättning",
"hälsomat",
"organist",
"vitaminer",
"hälsokost",
"köttersättning",
"vegetarian",
"hälsokostbutik"
],
"shop/hearing_aids":[
"hörselskada",
"hörapparater",
"Hörapparater",
"hörselskadade",
"hörsel",
"hörhjälpmedel"
],
"shop/herbalist":[
"läkande örter",
"örter",
"medicinalväxter",
"Medicinalväxter"
],
"shop/hifi":[
"ljudåtergivning",
"hifi",
"förstärkare",
"stereoanläggning",
"högtalare",
"HiFi-butik",
"ljudanläggning",
"stereo",
"hifi-butik",
"audio",
"video",
"ljud"
],
"shop/hobby":[
"hobbyaffär",
"Hobbyaffär",
"manga",
"model",
"modelljärnväg",
"modellflyg",
"hobby",
"modellbygge"
],
"shop/household_linen":[
"servetter",
"sängtextilier",
"linne",
"näsdukar",
"gardiner",
"bäddning",
"affär för hushållstextilier",
"Affär för hushållstextilier",
"filtar",
"handdukar",
"påslakan",
"överkast",
"textilier",
"dukar",
"lakan",
"örngott",
"hushållstextilier",
"kläder"
],
"shop/houseware":[
"porslin",
"hem",
"köksredskap",
"hushåll",
"husgeråd",
"bestick",
"prydnadsföremål",
"Husgeråd"
],
"shop/hunting":[
"jakt",
"Jaktbutik",
"jaktbutik",
"jaktaffär",
"jaktutrustning",
"jaktgevär",
"jaktvapen"
],
"shop/interior_decoration":[
"Inredningsaffär",
"inredning",
"inredningsaffär",
"dekoration"
],
"shop/jewelry":[
"pärla",
"ringar",
"armband",
"Juvelerare",
"ring",
"klockor",
"juvelerare",
"pärlor",
"halsband",
"diamant",
"smycken",
"guld",
"klocka",
"örhängen",
"silver",
"örhänge"
],
"shop/kiosk":[
"glass",
"gatukök",
"läsk",
"dryck",
"tobak",
"tidningar",
"snus",
"snabbmat",
"butik",
"godis",
"korv",
"cigaretter",
"Kiosk",
"kiosk"
],
"shop/kitchen":[
"kök",
"köksinredning",
"bänkskivor",
"köksskåp",
"skåpluckor",
"Köksinredning"
],
"shop/laundry":[
"Tvättinrättning",
"tvättomat",
"tvättstuga",
"tvättemat",
"tvättinrättning",
"tvättautomat",
"tvätt",
"tvätteri"
],
"shop/laundry/self_service":[
"tvättinrättning med självbetjäning",
"tvättomat",
"tvättstuga",
"tvättemat",
"tvättinrättning",
"tvättautomat",
"tvätt",
"Tvättinrättning med självbetjäning",
"tvätteri",
"mynttvätt"
],
"shop/leather":[
"läder",
"läderjackor",
"läderkläder",
"Läderaffär",
"läderaffär"
],
"shop/lighting":[
"belysningsbutik",
"led",
"belysning",
"lampor",
"glödlampor",
"Belysningsbutik"
],
"shop/locksmith":[
"låssmed",
"dyrkning",
"nyckel",
"nyckelkopiering",
"Låssmed",
"lås",
"låsinstallation",
"nyckeltillverkning",
"låsdyrkning"
],
"shop/lottery":[
"lottförsäljningen",
"bingospel",
"lottstånd",
"Lotteri",
"lotteri",
"hasardspel",
"hasard",
"lottdragning",
"tombola"
],
"shop/mall":[
"Köpcenter",
"shoppingcentrum",
"köpcentrum",
"köpcenter",
"shoppingcenter",
"varuhus",
"affärshus"
],
"shop/massage":[
"massagebehandling",
"thaimassage",
"Massage",
"massage"
],
"shop/medical_supply":[
"medicinsk utrustning",
"rullstol",
"blodtrycksmätare",
"kryckor",
"ortopedteknik",
"glucometer",
"hjälpmedel",
"ledstöd",
"glukometer",
"träningsbollar",
"Medicinsk utrustning",
"bandage"
],
"shop/military_surplus":[
"armé",
"krigsöverskott",
"affär med militäröverskott",
"vapen",
"militärutrustning",
"militärt överskott",
"militärkläder",
"överskottslagret",
"arméöverskott",
"marinöverskott",
"militäröverskott",
"Affär med militäröverskott",
"militär"
],
"shop/mobile_phone":[
"mobiltelefon",
"Mobiltelefoner",
"mobiltelefoni",
"telefon",
"mobiltelefoner",
"telefonbutik",
"mobiltelefonbutik"
],
"shop/model":[
"modellbyggnad",
"Affär för byggmodeller",
"modellbutik",
"skalmodeller",
"modellfigurer",
"modellpaket",
"modellbåtar",
"modellflyg",
"hobby",
"modellbygge"
],
"shop/money_lender":[
"utlåningsinstitution",
"telefonlån",
"mikrolån",
"pantbank",
"Långivare",
"utlåning",
"långivare"
],
"shop/motorcycle":[
"motorcykelbutik",
"motorcyklar",
"Återförsäljare av motorcyklar",
"motorcykeltillbehör",
"motorcykel",
"motorcykelåterförsäljare"
],
"shop/motorcycle_repair":[
"motorcykel",
"Motorcykelverkstad",
"motorcykelverkstad",
"motorcykelservice",
"verkstad",
"reparation",
"mopedverkstad",
"motorcykelreparatör",
"motorcyklar",
"service",
"cykel",
"moped",
"reparatör"
],
"shop/music":[
"cd",
"Musikaffär",
"kassett",
"lp",
"musikbutik",
"skivaffär",
"cd-affär",
"musikaffär",
"vinyl",
"skivbutik"
],
"shop/musical_instrument":[
"musikinstrument",
"noter",
"instrument",
"Musikinstrument"
],
"shop/newsagent":[
"pressbyrå",
"tidskrifter",
"tidningsaffär",
"Tidningsaffär",
"pressbyrån",
"tidningar",
"kiosk",
"magasin",
"tidningsställ",
"tidningskiosk"
],
"shop/nutrition_supplements":[
"viktminskning",
"hälsokost",
"hälsoörter",
"Hälsokost",
"hälsoprodukter",
"hälsa",
"mineraler",
"vitaminer"
],
"shop/optician":[
"glasögon",
"ögon",
"optiker",
"synundersökning",
"linser",
"Optiker"
],
"shop/outdoor":[
"tält",
"camping",
"klätterutrustning",
"vandring",
"klättring",
"vandringsutrustning",
"uteliv",
"friluftsaffär",
"campingutrustning",
"friluftsliv",
"Friluftsaffär"
],
"shop/outpost":[
"utlämning av online-beställningar",
"paketutlämning",
"online",
"posten",
"Utlämning av online-beställningar",
"internet",
"utlämning",
"paket"
],
"shop/paint":[
"färg",
"färgbutik",
"målarfärg",
"Färgbutik",
"målning"
],
"shop/party":[
"partyutrustning",
"partybutik",
"utklädning",
"kallasdekoration",
"festival",
"kallas",
"festivalutrustning",
"Partybutik",
"fest",
"engångstallrikar",
"festutrustning",
"ballonger",
"småpresenter",
"engångsbestick",
"dräkter",
"kallasutrustning",
"serpentiner",
"party",
"engångsglas",
"dekoration"
],
"shop/pastry":[
"kondis",
"kaffeservering",
"servering",
"fik",
"sockerbagare",
"kafé",
"konditori",
"café",
"finbageri",
"sockerbageri",
"cafe",
"bageri",
"Konditori"
],
"shop/pawnbroker":[
"pant",
"Pantbank",
"pantbelåning",
"pantbanken",
"pantbank",
"pantlånekontor",
"varubelåning"
],
"shop/perfumery":[
"parfymeri",
"Parfymbutik",
"parfym",
"parfymbutik",
"smink",
"kosmetika"
],
"shop/pet":[
"katter",
"katt",
"Djurbutik",
"hundar",
"djurmat",
"djuraffär",
"djur",
"akvarium",
"hund",
"fisk",
"djurburar",
"husdjur",
"djurtillbehör"
],
"shop/pet_grooming":[
"hund",
"pälsvård för husdjur",
"pälsvård",
"hundvård",
"trimning",
"husdjur",
"Pälsvård för husdjur"
],
"shop/photo":[
"fotoaffär",
"framkallning",
"kameratillbehör",
"fotokamera",
"video",
"film",
"konvertering",
"bild",
"fotografi",
"foto",
"kameror",
"Fotoaffär",
"filmkamera",
"fotoredigering",
"kamera",
"ram"
],
"shop/pottery":[
"keramikaffär",
"krukor",
"vaser",
"Keramikaffär",
"keramik"
],
"shop/printer_ink":[
"butik för skrivarbläck",
"skrivare",
"faxbläck",
"toner",
"kopiator",
"skrivarbläck",
"skrivartoner",
"Butik för skrivarbläck",
"bläck",
"fax",
"kopieringsbläck"
],
"shop/psychic":[
"seare",
"Medium / Psykisk",
"parapsykologi",
"spåman",
"ande",
"klärvoajans",
"tarotkort",
"ockult",
"medium",
"spådom",
"klärvoajant",
"synsk",
"spiritist",
"spåkvinna",
"kristallkula",
"sierska",
"spådam",
"tarot",
"astrologi",
"siare"
],
"shop/pyrotechnics":[
"Fyrverkerier",
"tomtebloss",
"raketer",
"smällare",
"fyrverkerier",
"pyroteknik",
"nyårsraketer"
],
"shop/radiotechnics":[
"elektronikbutik",
"radiotillbehör",
"radiobutik",
"elektronik",
"elektronikkomponenter",
"Radio/Elektronikbutik",
"radio"
],
"shop/religion":[
"religiös",
"biblar",
"kyrkobutik",
"psalmböcker",
"Religiös butik",
"religion"
],
"shop/rental":[
"hyra",
"hyrbutik",
"låna",
"Hyrbutik",
"uthyrning"
],
"shop/repair":[
"reparera",
"renovera",
"trasig",
"reparatör",
"Reparatör",
"laga",
"verkstad"
],
"shop/scuba_diving":[
"Dykarbutik",
"dykning",
"dykarbutik",
"dykutrustning"
],
"shop/seafood":[
"hummer",
"räkor",
"fisk",
"ostron",
"bläckfisk",
"fiskaffär",
"krabba",
"skaldjur",
"fiskhandlare",
"musslor",
"Fiskaffär"
],
"shop/second_hand":[
"loppis",
"Second hand",
"loppmarknad",
"second hand",
"secondhand"
],
"shop/sewing":[
"symaskin",
"tyg",
"sy",
"garn",
"Sybutik",
"nå",
"sybutik. sömnadsbutik",
"tråd",
"sömnad"
],
"shop/shoe_repair":[
"skoreparation",
"skoreparatör",
"skomakare",
"skor",
"Skomakare"
],
"shop/shoes":[
"Skoaffär",
"skoaffär",
"skobutik",
"skor"
],
"shop/spices":[
"chili",
"wasabi",
"salt",
"peppar",
"örter",
"gurkmeja",
"Affär för kryddor",
"curry",
"kryddor",
"kanel",
"affär för kryddor",
"saffran",
"kryddbutik",
"ingefära"
],
"shop/sports":[
"sportutrustning",
"träningsutrustning",
"träningskläder",
"sportkläder",
"löpskor",
"träningsskor",
"Sportaffär",
"sportaffär"
],
"shop/stationery":[
"grattiskort",
"papper",
"kort",
"kuvert",
"kontorsmaterial",
"pennor",
"anteckningsböcker",
"pappersvaror",
"pappershandel",
"Pappershandel"
],
"shop/storage_rental":[
"förråd",
"långtidslager",
"förrådsutrymme",
"bilförvaring",
"hyrlager",
"magasinera",
"förvaring",
"husvagnsförvaring",
"Hyrlager",
"båtförvaring",
"säsongsförvaring",
"vinterförvaring",
"magasinering",
"möbelförvaring"
],
"shop/supermarket":[
"supermarket",
"Mataffär",
"mat",
"snabbköp",
"självbetjäningsbutik",
"affär",
"livsmedelsbutik",
"mataffär",
"självköp",
"dagligvarubutik",
"livsmedel"
],
"shop/supermarket/organic":[
"supermarket",
"mat",
"snabbköp",
"Organisk mataffär",
"naturligt",
"naturlig mat",
"organisk mataffär",
"organisk mat",
"mataffär",
"organiskt"
],
"shop/swimming_pool":[
"basäng",
"poolinstallation",
"Butik för pooltillbehör",
"pool",
"poolbutik",
"pooltillbehörsbutik",
"poolservice",
"poolunderhåll",
"poolinstallationsbutik",
"jacussy",
"poolbutikleveransbutik´",
"badtunna",
"poolunderhållsbutik",
"poolutrustningsbutik"
],
"shop/tailor":[
"kostym",
"skräddare",
"klänning",
"kläder",
"Skräddare"
],
"shop/tattoo":[
"Tatueringsstudio",
"tatuera",
"tatuering",
"tatueringssalong",
"tatuerare",
"tatueringsstudio"
],
"shop/tea":[
"the",
"te",
"teblad",
"thé",
"örtte",
"Te-butik",
"påste"
],
"shop/telecommunication":[
"talkommunikation",
"röst",
"telekombutik",
"telefon",
"isp",
"internetleverantör",
"Telekombutik",
"tele",
"nätverk",
"internet",
"kommunikation"
],
"shop/ticket":[
"biljettlucka",
"biljettkassa",
"biljettkontor",
"biljetter",
"biljettsäljare",
"Biljettförsäljning",
"biljettförsäljning",
"biljettåterförsäljare"
],
"shop/tiles":[
"klinker",
"kakelplatta",
"plattsättare",
"plattor",
"Kakelbutik",
"kakelbutik",
"kakel"
],
"shop/tobacco":[
"tobaksbutik",
"pipor",
"cigarett",
"röktillbehör",
"tobak",
"cigarr",
"Tobaksbutik",
"cigaretter",
"snus",
"rökning",
"pipa",
"cigarrer"
],
"shop/tool_hire":[
"Verktygsuthyrning",
"byggverktyg",
"verktygsuthyrning",
"uthyrning av verktyg",
"hyrning",
"verktyg",
"byggmaskiner",
"uthyrning"
],
"shop/toys":[
"leksaker",
"leksaksaffär",
"barnsaker",
"Leksaksaffär"
],
"shop/trade":[
"Proffshandel",
"granngården",
"trävaror",
"trähandel",
"fönster",
"kakel",
"vvs-specialist",
"jordbruksprodukter",
"proffshandel",
"proffsmarknad",
"vvs",
"jordbruk",
"brädor",
"byggmaterial",
"lantmannaföreningen",
"brädgård",
"byggnadsmaterial",
"proffs"
],
"shop/travel_agency":[
"charterflyg",
"charter",
"resebyrå",
"reseagent",
"biljettförsäljning",
"charterresa",
"Resebyrå"
],
"shop/trophy":[
"medaljer",
"affär för troféer",
"trofe",
"troféer",
"Affär för troféer",
"plackat",
"trofé",
"priser",
"utmärkelser",
"trofeer",
"belöningar",
"gravyrer",
"trofébutik"
],
"shop/tyres":[
"däckförsäljning",
"däckbyte",
"hjulbyte",
"fälgar",
"däck",
"fälg",
"hjul",
"hjulförsäljning",
"balansering",
"Däckfirma",
"däckfirma"
],
"shop/vacant":[
"Tom lokal"
],
"shop/vacuum_cleaner":[
"dammsugarbutik",
"dammsugaråterförsäljare",
"dammsugarpåsar",
"Dammsugarbutik",
"dammsugartillbehör",
"dammsugare"
],
"shop/variety_store":[
"överskott",
"Fyndbutik",
"lågprisbutik",
"fynd",
"fyndbutik",
"billigt",
"lågpris",
"överskottsaffär"
],
"shop/video":[
"vhs",
"filmbutik",
"filmförsäljning",
"dvd",
"videobutik",
"Videobutik",
"filmuthyrning"
],
"shop/video_games":[
"tvspel",
"tv-spel",
"TV-spel",
"konsolspel",
"spelkonsoler",
"datorspel",
"videospel",
"dataspel"
],
"shop/watches":[
"klockaffär",
"Klockaffär",
"klockbutik",
"klocka",
"klockor",
"uraffär",
"urbutik",
"ur"
],
"shop/water":[
"dricksvatten",
"Affär för dricksvatten",
"vatten"
],
"shop/water_sports":[
"simning",
"badkläder",
"Vattensport/simning",
"vattensport"
],
"shop/weapons":[
"ammunition",
"jakt",
"skjutvapen",
"vapen",
"kniv",
"knivar",
"pistol",
"vapenaffär",
"Vapenaffär"
],
"shop/wholesale":[
"grosshandel",
"grossistverksamhet",
"engros",
"mängdhandel",
"lagerklubb",
"grosist",
"grossistklubb",
"Grosistaffär",
"partihandel",
"grossistlager",
"grosistaffär"
],
"shop/wigs":[
"peruker",
"Affär för peruker",
"hårförlängning",
"löshår",
"tupé",
"affär för peruker"
],
"shop/window_blind":[
"spjälgardin",
"spjäljalusi",
"Persienner",
"markis",
"persienner",
"jalusi",
"rullgardin"
],
"shop/wine":[
"vinaffär",
"systemet",
"systembolaget",
"vin",
"vinförsäljning",
"Vinaffär"
],
"telecom":[
"Telekomobjekt"
],
"telecom/data_center":[
"datasystem",
"datorcenter",
"datacenter",
"it",
"serverfarm",
"telekommunikation",
"serverhall",
"it-center",
"informationsteknologi",
"datorsystem",
"Datacenter",
"serverrum",
"molnet",
"datalagring"
],
"telecom/exchange":[
"telefonstation",
"Telefonstation",
"telefonväxel",
"telekommunikation"
],
"tourism":[
"Turistobjekt"
],
"tourism/alpine_hut":[
"fjällstuga",
"Fjällstation",
"fjällstation"
],
"tourism/apartment":[
"turist",
"hotell",
"turistlägenhet",
"andelslägenhet",
"gästlägenhet",
"condo",
"Turistlägenhet",
"lägenhetshotell",
"lägenhet"
],
"tourism/aquarium":[
"akvarium",
"fisk",
"Akvarium",
"hav",
"vatten"
],
"tourism/artwork":[
"Publik konst",
"målning",
"konst",
"gatukonst",
"väggmålning",
"offentlig konst",
"publik konst",
"skulptur",
"staty"
],
"tourism/artwork/bust":[
"byst",
"Byst",
"figur",
"staty"
],
"tourism/artwork/graffiti":[
"klotter",
"spray",
"Graffiti",
"graffitikonst",
"kladd",
"sprayfärg",
"graffiti",
"gatukonst"
],
"tourism/artwork/installation":[
"konstinstallation",
"interaktiv konst",
"kultur",
"installation",
"modern konst",
"konst",
"Konstinstallation"
],
"tourism/artwork/mural":[
"fresco",
"mural",
"målning",
"Väggmålning",
"väggmålning"
],
"tourism/artwork/sculpture":[
"byst",
"Skulptur",
"monument",
"snideri",
"staty",
"skulptur",
"figur"
],
"tourism/artwork/statue":[
"Staty",
"byst",
"monument",
"snideri",
"staty",
"skulptur",
"figur"
],
"tourism/attraction":[
"Turistattraktion",
"sevärdighet",
"turistattraktion",
"sevärdhet"
],
"tourism/camp_pitch":[
"tält",
"tältplats",
"camping",
"husvagn",
"Tältplats/husvagnsplats",
"husvagnsplats",
"campingplats"
],
"tourism/camp_site":[
"tält",
"campinganläggning",
"camping",
"husvagn",
"Campingplats",
"campingplats"
],
"tourism/camp_site/backcountry":[
"vildmark",
"enkel camping",
"Vildmarkscamping",
"primitiv camping",
"friluftscamping",
"naturcamping",
"informell camping",
"vildmarkscamping",
"campingplats"
],
"tourism/camp_site/group_only":[
"Gruppcampingplats",
"gruppcampingplats",
"campingplats för grupp",
"lägerplats",
"campingplats",
"scoutcamping",
"ungdomscamping"
],
"tourism/caravan_site":[
"camping",
"husvagnscamping",
"husbilscamping",
"ställplats",
"Ställplats",
"campingplats",
"fricamping"
],
"tourism/chalet":[
"helgboende",
"camping",
"stuga",
"sommarstuga",
"Stuga",
"helg",
"campingstuga",
"semester",
"semesterboende",
"semesterstuga",
"ledighet"
],
"tourism/gallery":[
"konstaffär",
"Konstgalleri",
"konstverk",
"tavlor",
"kulturer",
"konst",
"konsthandlare",
"konstgalleri",
"galleri",
"statyer",
"konstutställning"
],
"tourism/guest_house":[
"b&d",
"vandrarhem",
"gästhus",
"logi",
"bed & breakfast",
"övernattningsställe",
"pensionat",
"Gästhus"
],
"tourism/hostel":[
"Vandrarhem",
"vandrarhem",
"övernattningsställe"
],
"tourism/hotel":[
"hotell",
"värdshus",
"Hotell",
"hotellanläggning"
],
"tourism/information":[
"infokarta",
"karta",
"informationskarta",
"information",
"Information",
"turistkontor",
"informationstavla",
"informationskällan",
"turistbyråer"
],
"tourism/information/board":[
"turistinformation",
"avgång*",
"kollektivtrafik",
"fakta",
"karta",
"Informationstavla",
"information",
"historisk information",
"informationstavla"
],
"tourism/information/board/welcome_sign":[
"välkomstskylt",
"välkomna",
"välkommen",
"Välkomstskylt",
"skylt"
],
"tourism/information/guidepost":[
"guidepost",
"stigvisning",
"Vägvisare",
"vandringsskyllt",
"vägvisare",
"vägmärke"
],
"tourism/information/map":[
"*karta",
"cykelkarta",
"Karta",
"karta",
"navigering",
"information",
"stadskarta",
"vägkarta",
"informationstavla",
"industrikarta"
],
"tourism/information/office":[
"turist",
"Turistbyrå",
"turistinformationscenter",
"informationskontor",
"turism",
"besöksinformationscenter",
"turistkontor",
"reseguide",
"turistinformation",
"turistbyrå",
"resebyrå",
"besökscenter",
"välkomstcenter"
],
"tourism/information/route_marker":[
"skidled",
"ridled",
"stigmarkör",
"vandring",
"ledmarkör",
"vägmarkör",
"skoterled",
"stig",
"led",
"ruttflagga",
"ruttmarkör",
"stenhög",
"Spårmarkör",
"rutt",
"vandringsled",
"spår",
"spårmarkör"
],
"tourism/information/terminal":[
"informationsterminal",
"infokarta",
"turistbyrå",
"turistkartor",
"Informationsterminal",
"informationskälla",
"karta",
"informationskarta",
"information",
"terminal"
],
"tourism/motel":[
"motorhotell",
"motell",
"hotell",
"väghotell",
"Motel"
],
"tourism/museum":[
"samling",
"museibyggnad",
"historia",
"museum",
"vetenskap",
"utställning",
"konstsamling",
"Museum",
"historik",
"konst",
"arkeologi",
"galleri"
],
"tourism/museum/history":[
"diorama",
"historia",
"grund",
"historisk",
"utställning",
"Historiskt museum",
"hall",
"utställningar",
"artefakter",
"institution",
"museum",
"historiskt museum",
"stadsmuseum"
],
"tourism/picnic_site":[
"Picknickplats",
"picknickplats",
"camping",
"rastplats",
"utflykt",
"campingplats",
"picknick"
],
"tourism/theme_park":[
"nöjespark",
"temapark",
"åkattraktioner",
"nöjesplats",
"tivoli",
"nöjesfält",
"Nöjespark"
],
"tourism/trail_riding_station":[
"tur",
"ridstation",
"hästrastning",
"häststall",
"gästhus",
"ridningsstation",
"stall",
"turridningsstation",
"turridning",
"Turridningsstation",
"häst"
],
"tourism/viewpoint":[
"utsikt",
"vy",
"utsiktsplats",
"Utsiktspunkt"
],
"tourism/wilderness_hut":[
"hydda",
"vandring",
"ödestuga",
"stuga",
"skydd",
"koja",
"hajk",
"kyffe",
"övernattning",
"Stuga (för vandrare o.d.)",
"vildmarksstuga",
"barack",
"fjällstuga",
"stuga (för vandrare o.d.)",
"fjällstation"
],
"tourism/zoo":[
"djurpark",
"zoo",
"Zoo",
"zoologisk trädgård"
],
"tourism/zoo/petting":[
"barn-zoo",
"barn",
"mini-zoo",
"djurpark",
"klappa",
"klapp-zoo",
"minidjurpark",
"barndjurpark",
"zoo",
"djur",
"lantgårdsdjur",
"Barn-zoo"
],
"tourism/zoo/safari":[
"Safaridjurpark",
"safari",
"genomkörningsdjurpark",
"safaridjurpark",
"djurpark",
"zoo",
"safaripark"
],
"tourism/zoo/wildlife":[
"vilddjurspark",
"Vilddjurspark",
"djurpark",
"inhemska djur",
"vilddjur",
"zoo"
],
"traffic_calming":[
"långsam",
"hastighet",
"fartgupp",
"* fart*",
"farthinder",
"gupp",
"trafikhinder",
"säkerhet",
"Farthinder"
],
"traffic_calming/bump":[
"bula",
"Fartbula (kort gupp)",
"fartbula",
"bump",
"fartgupp",
"vägbula",
"farthinder",
"gupp"
],
"traffic_calming/chicane":[
"sidoförskjutning",
"trafikchikan",
"långsam",
"hastighet",
"* fart*",
"farthinder",
"Sidoförskjutning (chikan)",
"kurvor",
"chikan",
"slalom",
"trafikhinder",
"säkerhet"
],
"traffic_calming/choker":[
"lins",
"choker",
"Avsmalning",
"avsmalning",
"långsam",
"hastighet",
"* fart*",
"farthinder",
"trafikhinder",
"säkerhet",
"timglas"
],
"traffic_calming/cushion":[
"lins",
"vägkudde",
"långsam",
"hastighet",
"fartgupp",
"* fart*",
"farthinder",
"Vägkudde",
"trafikhinder",
"gupp",
"säkerhet",
"timglas"
],
"traffic_calming/dip":[
"långsam",
"hastighet",
"fartgupp",
"grop",
"* fart*",
"farthinder",
"trafikhinder",
"Grop",
"säkerhet",
"försänkning"
],
"traffic_calming/hump":[
"normalt fartgupp",
"cirkulärt gupp",
"wattgupp",
"wattska guppet",
"gp-gupp",
"fartpuckel",
"puckel",
"fartgupp",
"farthinder",
"Normalt fartgupp",
"standardgupp",
"gupp"
],
"traffic_calming/island":[
"cirkulation",
"långsam",
"hastighet",
"cirkel",
"sidorefug",
"refug",
"mittrefug",
"trafikö",
"ö",
"Refug",
"cirkulationsplats",
"* fart*",
"farthinder",
"trafikhinder",
"säkerhet",
"rondell"
],
"traffic_calming/rumble_strip":[
"pennsylvaniaräfflor",
"Bullerräfflor",
"bullerräfflor"
],
"traffic_calming/table":[
"fartgupp (långt)",
"Fartgupp (långt)",
"fartgupp",
"farthinder",
"platågupp",
"långt fartgupp",
"gupp"
],
"traffic_sign":[
"Vägmärke",
"trafikskyllt",
"trafikmärke",
"skyllt",
"vägskyllt",
"vägmärke",
"vägvisare"
],
"traffic_sign/city_limit":[
"Skyllt för tättbebyggt område",
"trafikskyllt",
"tättbebyggt område",
"skyllt",
"stadsgräns",
"ort",
"stad",
"tätort",
"trafikmärke",
"gräns",
"vägskyllt",
"vägmärke",
"vägvisare"
],
"traffic_sign/maxspeed":[
"trafikskyllt",
"hastighetsskylt",
"skyllt",
"hastighet",
"fart",
"maxhastighet",
"trafikmärke",
"maxfart",
"Hastighetsskylt",
"vägskyllt",
"hastighetsbegränsning",
"vägmärke",
"vägvisare"
],
"type/boundary":[
"gränslinje",
"Gräns",
"administrativ gräns",
"gräns"
],
"type/boundary/administrative":[
"stat",
"Administrativ gräns",
"administrativ gräns",
"administrativ enhet",
"gräns",
"territorium"
],
"type/connectivity":[
"Filkoppling",
"filer",
"sammankoppling av filer",
"filkoppling",
"vägfil",
"anslutning",
"filbyte"
],
"type/destination_sign":[
"vägvisning",
"vägskylt",
"Destinationsskylt",
"destination",
"destinationsskylt",
"skylt",
"vägvisare"
],
"type/enforcement":[
"fartkontroll",
"fartkamera",
"hastighetskamera",
"Trafiksäkerhetsutrustning",
"trafiksäkerhet",
"övervakning",
"hastighetskontroll",
"trafiksäkerhetsutrustning"
],
"type/enforcement/maxspeed":[
"fartkamera",
"hastighetskamera",
"fartkontroll",
"fart",
"radar",
"trafiksäkerhetskamera",
"trafiksäkerhet",
"Fartkamera",
"övervakning",
"hastighetskontroll",
"hastighet",
"trafiksäkerhetsutrustning"
],
"type/multipolygon":[
"Multipolygon"
],
"type/public_transport/stop_area_group":[
"Grupp av stopp för kollektivtrafik",
"kollektivtrafik",
"hållplats",
"bytespunkt",
"transit",
"byte",
"station",
"knutpunkt",
"resecenter",
"terminal",
"linjetrafik",
"transport"
],
"type/restriction":[
"restriktion",
"begränsning",
"inskränkning",
"förbehåll",
"Restriktion"
],
"type/restriction/no_left_turn":[
"ingen vänstersväng",
"Ingen vänstersväng",
"sväng ej vänster"
],
"type/restriction/no_right_turn":[
"ingen högersväng",
"ej högersväng",
"sväng ej höger",
"Ingen högersväng"
],
"type/restriction/no_straight_on":[
"ej rakt fram",
"Ej rakt fram",
"fortsätt ej framåt"
],
"type/restriction/no_u_turn":[
"ingen u-sväng",
"får ej vända",
"Ingen U-sväng"
],
"type/restriction/only_left_turn":[
"enbart vänstersväng",
"vänster",
"Enbart vänstersväng",
"vänstersväng"
],
"type/restriction/only_right_turn":[
"Enbart högersväng",
"högersväng",
"höger",
"enbart högersväng"
],
"type/restriction/only_straight_on":[
"Enbart rakt fram",
"fortsätt framåt",
"får ej svänga",
"enbart rakt fram"
],
"type/restriction/only_u_turn":[
"u-sväng",
"måste vända",
"Enbart U-sväng",
"enbart u-sväng"
],
"type/route":[
"Rutt",
"rutt",
"färdled",
"färdväg"
],
"type/route/aerialway":[
"rutt för linbana",
"linbanerutt",
"linbana",
"Linbanerutt"
],
"type/route/bicycle":[
"cykelled",
"cykelförbindelse",
"cykelnät",
"Cykelrutt",
"cykelrutt"
],
"type/route/bus":[
"busslinje",
"bussväg",
"Busslinje",
"bussrutt",
"bussled"
],
"type/route/detour":[
"Alternativ rutt",
"alternativ rutt",
"omväg",
"alternativ väg"
],
"type/route/ferry":[
"båtrutt",
"båtlinjetrafik",
"Färjerutt",
"färjerutt"
],
"type/route/foot":[
"Vandringsled",
"gångled",
"vandring",
"gång",
"vandringsled",
"gångrutt",
"stig",
"vandringsrutt"
],
"type/route/hiking":[
"Vandringsled",
"vandringsled",
"stig",
"vandringsrutt"
],
"type/route/horse":[
"rida",
"ridled",
"ridturism",
"ridning",
"hästled",
"häst",
"ridväg",
"hästsport",
"hästväg",
"långfärdsridning",
"ridrutt",
"Ridled",
"ridetapp",
"hästrutt"
],
"type/route/light_rail":[
"tågrutt",
"smalspårig järnväg",
"rutt för snabbspårväg",
"järnvägsförbindelse",
"stadsbana",
"järnvägsrutt",
"rutt på smalspårig järnväg",
"snabbspårväg",
"smalspår",
"Rutt på snabbspårväg / stadsbana",
"tågnät",
"rutt för stadsbana",
"järnväg"
],
"type/route/monorail":[
"Monorailrutt",
"kollektivtrafik",
"enskensbana",
"linjetrafik",
"transport",
"balkbana",
"spår",
"räls",
"monorail"
],
"type/route/mtb":[
"enduro",
"mountainbikerutt",
"Mountainbikerutt",
"terrängcykling",
"freeride",
"trail ridning",
"mtb",
"mountainbike",
"utförsåkning"
],
"type/route/pipeline":[
"pipeline",
"oljeledning",
"vattenledning",
"avloppsledning",
"rörledningsrutt",
"rörledning",
"Rörledningsrutt"
],
"type/route/piste":[
"längdskidspår",
"pistspår",
"Pist/skidrutt",
"skidor",
"skidtur",
"snöpark",
"skidbacke",
"utförsåkning",
"pist",
"skridskorutt",
"skidrutt",
"slädspår",
"längdskidåkning",
"slalombacke",
"skidspår",
"skidbana",
"skridskospår",
"skridskobana"
],
"type/route/power":[
"kraftledningsrutt",
"kraftledning",
"elnät",
"Kraftledningsrutt",
"elförsörjning"
],
"type/route/road":[
"Vägrutt",
"vägförbindelse",
"vägnät",
"vägrutt"
],
"type/route/subway":[
"Tunnelbanerutt",
"tunnelbanerutt",
"tunnelbana"
],
"type/route/train":[
"tågrutt",
"tågnät",
"järnvägsförbindelse",
"Tågrutt",
"järnväg",
"järnvägsrutt"
],
"type/route/tram":[
"spårvagnsrutt",
"spårvagnsnät",
"Spårvagnsrutt",
"spårvagn",
"spårvagnsförbindelse",
"spårvagnsräls"
],
"type/route/trolleybus":[
"Trådbussrutt",
"trådbuss",
"trådbussrutt",
"kollektivtrafik",
"spårlös",
"bussrutt",
"transit",
"spårvagn",
"transport",
"buss",
"vag"
],
"type/route_master":[
"huvudrutt",
"huvudförbindelse",
"huvudväg",
"Huvudrutt"
],
"type/site":[
"anläggning",
"läge",
"plats",
"ställe",
"Plats"
],
"type/waterway":[
"vattenväg",
"vattendrag",
"Vattendrag",
"vattenflöde"
],
"waterway":[
"Vattenvägobjekt"
],
"waterway/boatyard":[
"båtvarv",
"båtställplats",
"varv",
"Båtvarv",
"uppläggningsplats",
"vinterförvaring"
],
"waterway/canal":[
"vattenväg",
"kanal",
"vattenled",
"Kanal"
],
"waterway/canal/lock":[
"ränna",
"slusskammare",
"slussbassäng",
"vattenlås",
"Sluss",
"kanalsluss",
"sluss"
],
"waterway/dam":[
"fördämning",
"vattensamling",
"damm",
"reservoar",
"Fördämning"
],
"waterway/ditch":[
"dike",
"fåra",
"Dike"
],
"waterway/dock":[
"båtdocka",
"båtvarv",
"fartygsvarv",
"Våt- / Torrdocka",
"varv",
"torrdocka",
"docka",
"lastdocka",
"våtdocka",
"fartygsdocka"
],
"waterway/drain":[
"dagvattenavrinning",
"dagvatten",
"Dränering",
"dränering",
"avrinning"
],
"waterway/fish_pass":[
"fisklås",
"fiskväg",
"ålstege",
"fisksteg",
"fisktrappa",
"fiskpassage",
"Fisktrappa",
"fiskstege",
"fiskvandring",
"ålpassering"
],
"waterway/fuel":[
"sjömack",
"båtmack",
"tankstation båtbensninmack",
"bränslestation",
"båtmensinstation",
"Sjömack"
],
"waterway/lock_gate":[
"slussport",
"kanal",
"Slussport",
"sluss"
],
"waterway/milestone":[
"Milsten vid vattendrag",
"kilometertavla",
"kilometerpåle",
"sjöfart",
"milsten",
"referenstavla",
"milsten vid vattendrag",
"kilometerstolpe",
"avståndsmärke"
],
"waterway/river":[
"vattendrag",
"ström",
"jokk",
"å",
"fors",
"Flod",
"flod",
"älv"
],
"waterway/riverbank":[
"Flodbank"
],
"waterway/sanitary_dump_station":[
"tömningsplats",
"båtlatrin",
"gråvatten",
"båtsanitet",
"gråvattentömning",
"Marin latrintömning",
"sanitet",
"latrintömning",
"vattenfarkoster",
"cdp",
"båttömnig",
"båt",
"sanitära",
"marin latrintömning",
"ctdp",
"kemisk toalett",
"toalettömning",
"pumpa ut",
"utpumpning",
"dumpstation",
"elsan",
"campingtoalett"
],
"waterway/stream":[
"dike",
"biflod",
"vattendrag",
"flöde",
"ström",
"bäck",
"biflöde",
"flod",
"Bäck",
"rännil"
],
"waterway/stream_intermittent":[
"Periodiskt vattendrag",
"bäck",
"periodiskt",
"arroyo",
"dagvatten",
"biflöde",
"tillfälligt",
"översvämning",
"dike",
"vattendrag",
"tillfälligt vattendrag",
"dränering",
"periodiskt vattendrag",
"avrinning",
"rännil"
],
"waterway/tidal_channel":[
"vattenväg",
"tidvattenbäck",
"tidvatten",
"Tidvattenskanal",
"kust",
"salt kärr",
"tidvattenskanal",
"tidvatteninlopp",
"marin"
],
"waterway/water_point":[
"dricksvatten för båt",
"dricksvatten",
"Dricksvatten för båt",
"vattenpåfyllning",
"vattentank"
],
"waterway/waterfall":[
"Vattenfall",
"fall",
"vattenfall",
"fors"
],
"waterway/weir":[
"fördämning",
"vattensamling",
"damm",
"reservoar",
"Damm"
]
}
