{
"address":[
"postadress",
"postnummer",
"husnummer",
"Adress",
"destination",
"gatuadress",
"postort"
],
"advertising/billboard":[
"affischtavla",
"reklamskylt",
"reklamtavla",
"affisch",
"reklam",
"Annonstavla"
],
"advertising/column":[
"annonstavla",
"reklamplats",
"Reklampelare",
"annons",
"affisch",
"reklam",
"affischpelare",
"reklampelare",
"billboard",
"marknadsföring",
"annonspelare",
"annonsering"
],
"aerialway":[
"Linbana"
],
"aerialway/cable_car":[
"Kabinbana",
"linbana",
"pendelbana"
],
"aerialway/chair_lift":[
"lift",
"linbana",
"Expresslift",
"Stollift",
"stolslift",
"skidlift"
],
"aerialway/drag_lift":[
"Släplift",
"Draglift",
"lift",
"linbana",
"skidlift"
],
"aerialway/gondola":[
"Gondolbana",
"lift",
"linbana",
"Gondol",
"skidlift"
],
"aerialway/goods":[
"gruvlift",
"transportbana",
"varor",
"gods",
"varulift",
"linbana",
"transport",
"industrilift",
"Transportlift",
"transportlinbana",
"lift",
"industri",
"Transportlinbana"
],
"aerialway/magic_carpet":[
"skidliften",
"släplift",
"lift",
"Rullband",
"magisk matta"
],
"aerialway/mixed_lift":[
"Hybridlift (Telemixlift)",
"stollift",
"expresslift",
"Telemixlift",
"gondol",
"lift",
"linbana",
"skidlift",
"stolslift",
"hybridlift",
"gondolbana"
],
"aerialway/platter":[
"tallrikslift",
"släplift",
"lift",
"knapp",
"linbana",
"tallrik",
"Knapplift",
"skidlift"
],
"aerialway/pylon":[
"pylon",
"stolpe",
"Linbanestolpe",
"stötta",
"pelare"
],
"aerialway/rope_tow":[
"släplift",
"lift",
"linbana",
"skidlift",
"Replift"
],
"aerialway/station":[
"Linbanestation"
],
"aerialway/t-bar":[
"Ankarlift",
"släplift",
"T-lift",
"lift",
"linbana",
"skidlift",
"T-bygellift"
],
"aeroway":[
"Flygtrafik"
],
"aeroway/aerodrome":[
"flyghamn",
"flyg",
"flygplats",
"aerodrom",
"Flygplats",
"lufthamn",
"flygfält",
"flygplan",
"landningsplats"
],
"aeroway/apron":[
"flygparkering",
"Flygplansparkering",
"parkering av flygplan",
"apron",
"Parkering av flygplan (Apron)",
"parkering av plan",
"flygplansplatta",
"flygplatsplatta"
],
"aeroway/gate":[
"flyggate",
"flygplatsgate",
"Gate"
],
"aeroway/hangar":[
"Hangar",
"flygverkstad",
"flygplansgarage",
"flyggarage",
"garage för flygplan",
"flygplanshall"
],
"aeroway/helipad":[
"Helipad",
"Helikopterplatta",
"helikopter"
],
"aeroway/runway":[
"Start- och landningsbana",
"landningsbana",
"Startbana",
"landa",
"landning",
"rullbana"
],
"aeroway/taxiway":[
"flygplansväg",
"transportbana",
"Taxibana",
"transportsträcka"
],
"aeroway/terminal":[
"flygplats",
"Flygterminal",
"Flygplatsterminal",
"flygterminal",
"terminal",
"avgångshall",
"ankomsthall"
],
"allotments/plot":[
"odlingslott",
"lott",
"koloniträdgård",
"koloniområde",
"Kolonilott",
"koloni",
"täppa"
],
"amenity":[
"Facilitet"
],
"amenity/animal_boarding":[
"kattpensionat",
"katt",
"hundkollo",
"Djurhotell",
"katthotell",
"häst",
"Hundhotell",
"hund",
"Hundpensionat",
"inackordering",
"reptil",
"djurkollo",
"Djurpensionat",
"husdjur",
"kattkollo"
],
"amenity/animal_breeding":[
"katt",
"ko",
"tjur",
"kattunge",
"djurhållning",
"häst",
"avel",
"hund",
"reptil",
"valp",
"boskap",
"Djuruppfödning",
"djuravel",
"husdjur",
"Uppfödning",
"djuruppfödning"
],
"amenity/animal_shelter":[
"Djurhem",
"katthem",
"hemlös",
"katt",
"rovfågel",
"häst",
"vanvårdad",
"hund",
"reptil",
"omplacering",
"djuradoption",
"karantän",
"husdjur",
"omhändertagande",
"djurskydd"
],
"amenity/arts_centre":[
"kulturcenter",
"museum",
"kultur",
"tavlor",
"kulturhus",
"Konstcenter",
"konst"
],
"amenity/atm":[
"bankomat",
"minuten",
"otto",
"uttagsautomat",
"Uttagsautomat",
"atm",
"kontanter",
"pengar"
],
"amenity/bank":[
"kreditinrättning",
"investering",
"Bank",
"bankkontor",
"insättning",
"check",
"låneinstitut",
"bankvalv",
"besparing",
"penninginrättning",
"fonder",
"banklokal",
"kassa",
"penninganstalt"
],
"amenity/bar":[
"Bar",
"matställe",
"servering",
"saloon",
"öl",
"cocktailsalong",
"sprit",
"pub",
"krog"
],
"amenity/bbq":[
"bbq",
"Grill",
"eldning",
"eldstad",
"Barbecue",
"grillplats",
"Grillplats/Grill",
"eldplats",
"grillning"
],
"amenity/bench":[
"sits",
"bänk",
"sittmöbel",
"sittbräde",
"soffa",
"Bänk"
],
"amenity/bicycle_parking":[
"ställplats",
"cykel",
"Cykelparkering",
"cykelställ",
"Parkering"
],
"amenity/bicycle_rental":[
"Cykeluthyrning",
"lånecykel",
"cykellån",
"cykel",
"cykelleasing",
"hyrcykel"
],
"amenity/bicycle_repair_station":[
"Cykelreparation",
"kedjebrytare",
"Station för cykelreparation",
"cykel",
"tryckluft",
"cykelpump",
"pumpstation"
],
"amenity/biergarten":[
"ölträdgård",
"servering",
"trädgårdsbar",
"sprit",
"krog",
"utepub",
"utecafé",
"bar",
"Ölträdgård",
"Biergarten",
"utebar",
"öl",
"pub",
"trädgårdspub",
"uteservering",
"ölcafé"
],
"amenity/boat_rental":[
"båtleasing",
"lånebåt",
"Båtuthyrning",
"hyrbåt",
"båtlån"
],
"amenity/bureau_de_change":[
"resecheckar",
"valuta",
"pengaväxlare",
"Växlingskontor",
"pengaväxling",
"växling",
"pengar"
],
"amenity/bus_station":[
"Busstation / Bussterminal"
],
"amenity/cafe":[
"te",
"kondis",
"kaffeservering",
"servering",
"kaffestuga",
"kafeteria",
"fik",
"cafeteria",
"konditori",
"bistro",
"kaffe",
"Café"
],
"amenity/car_pooling":[
"lånebil",
"hyrbil",
"Bilpool"
],
"amenity/car_rental":[
"Biluthyrning",
"lånebil",
"hyrbil",
"billån",
"billeasing"
],
"amenity/car_sharing":[
"bildelning",
"Bilpool"
],
"amenity/car_wash":[
"biltvättanläggning",
"tvättgata",
"tvätt-tunnel",
"portaltvätt",
"Biltvätt"
],
"amenity/casino":[
"Tärning",
"spelsalong",
"Kasino",
"poker",
"spelklubb",
"spelhåla",
"spelrum",
"blackjack",
"kasino",
"spelhus",
"spel",
"Casino",
"roulette",
"kortspel",
"hasardspel"
],
"amenity/charging_station":[
"snabbladdning",
"eluttag",
"el",
"Laddstation",
"elbil"
],
"amenity/childcare":[
"lekgrupp",
"Förskola",
"Barnomsorg",
"daghem",
"Barnhem",
"Dagmamma",
"Dagis"
],
"amenity/cinema":[
"bioduk",
"Bio",
"Biografteater",
"film",
"Biograf",
"drive-in"
],
"amenity/clinic":[
"sjukvård",
"distriktssköterska",
"doktor",
"Klinik",
"vårdcentral",
"distriktsläkare",
"sjukhus",
"Vårdcentral",
"primärvård",
"läkare"
],
"amenity/clinic/abortion":[
"framkallat missfall",
"abort",
"Abortklinik",
"missfall",
"abortklinik",
"fosterfördrivning",
"avbrytande av havandeskap"
],
"amenity/clinic/fertility":[
"Insemination",
"Fertilitetscentrum",
"Fertilitet",
"barnlöshet",
"fortplantning",
"ägglossning",
"Äggfrys",
"spermie",
"spermadonation",
"befruktning",
"reproduktion",
"IVF",
"äggdonation",
"Fertilitetsklinik"
],
"amenity/clock":[
"väggur",
"urtavla",
"kyrkklocka",
"solur",
"Klocka",
"ur",
"väggklocka",
"tidur"
],
"amenity/college":[
"college",
"gymnasieområde",
"gymnasie",
"vidareutbildning",
"gymnasiumområde",
"Gymnasium",
"Collegeområde"
],
"amenity/community_centre":[
"folkets hus",
"bygdegård",
"Sockenstuga",
"Samlingslokal",
"folkets park",
"Hembygdsgård",
"byförening",
"festlokal",
"Byalag",
"bystuga",
"evenemang"
],
"amenity/compressed_air":[
"Tryckluft",
"pumpstation",
"komprimerad luft"
],
"amenity/courthouse":[
"lag",
"rätt",
"Domstol",
"juridik",
"ting",
"rättskipare",
"tribunal",
"instans",
"lagbok"
],
"amenity/coworking_space":[
"Dagkontor"
],
"amenity/crematorium":[
"begravning",
"Krematorium",
"kremering"
],
"amenity/dentist":[
"tänder",
"tanddoktor",
"odontolog",
"tandborstning",
"tand",
"Tandläkare",
"tandhygien",
"tandhygienist"
],
"amenity/dive_centre":[
"sportdykare",
"sportdykning",
"dykare",
"Dykcenter",
"scuba",
"dykning",
"grodman"
],
"amenity/doctors":[
"klinik",
"sjukvård",
"sjukvårdare",
"doktor",
"vårdcentral",
"sjukhus",
"läkare",
"Doktor",
"vårdinrättning"
],
"amenity/dojo":[
"Dojo",
"kampsport",
"budo",
"japan",
"japansk konst",
"Dojo / Akademi för kampsport",
"kampkonst",
"dojang",
"träningslokal"
],
"amenity/drinking_water":[
"Dricksvatten ",
"Dricksvatten",
"källa",
"fontän",
"vatten"
],
"amenity/driving_school":[
"bilskola",
"körkort",
"Trafikskola",
"uppkörning",
"lastbilskort",
"övningskörning",
"körskola"
],
"amenity/embassy":[
"legation",
"Ambassad",
"diplomatisk beskickning",
"utlandsrepresentation",
"beskickning",
"ambassad"
],
"amenity/fast_food":[
"skräpmat",
"Snabbmat",
"gatuköksmat",
"hämtmat",
"gatukök",
"restaurang",
"takeaway",
"bukfylla",
"junk-food"
],
"amenity/fast_food/burger":[
"mat",
"lunch",
"gatukök",
"restaurang",
"burgare",
"takeaway",
"bukfylla",
"junk-food",
"skräpmat",
"Snabbmat",
"gatuköksmat",
"hämtmat",
"äta",
"hamburgare",
"Snabbmat – Hamburgare",
"drive-in",
"grill"
],
"amenity/fast_food/chicken":[
"mat",
"Snabbmat – Kyckling",
"lunch",
"gatukök",
"restaurang",
"takeaway",
"bukfylla",
"junk-food",
"skräpmat",
"Snabbmat",
"gatuköksmat",
"hämtmat",
"äta",
"kyckling",
"drive-in",
"grill"
],
"amenity/fast_food/fish_and_chips":[
"mat",
"lunch",
"fisk och chips",
"gatukök",
"restaurang",
"Snabbmat – Fish & Chips",
"takeaway",
"bukfylla",
"junk-food",
"skräpmat",
"Snabbmat",
"gatuköksmat",
"hämtmat",
"äta",
"Fish and chips",
"Fish & chips",
"drive-in",
"grill"
],
"amenity/fast_food/kebab":[
"mat",
"lunch",
"gatukök",
"restaurang",
"takeaway",
"bukfylla",
"junk-food",
"skräpmat",
"Snabbmat",
"gatuköksmat",
"hämtmat",
"äta",
"kebab",
"Snabbmat – Kebab",
"drive-in",
"grill"
],
"amenity/fast_food/pizza":[
"mat",
"Snabbmat – Pizza",
"lunch",
"pan pizza",
"gatukök",
"restaurang",
"takeaway",
"bukfylla",
"junk-food",
"skräpmat",
"Snabbmat",
"gatuköksmat",
"hämtmat",
"äta",
"pizza",
"pizzeria",
"drive-in",
"grill"
],
"amenity/fast_food/sandwich":[
"lunch",
"smörgåsar",
"macka",
"bargetter",
"Snabbmat – Smörgås",
"skräpmat",
"Snabbmat",
"gatuköksmat",
"hämtmat",
"äta",
"smörgås",
"baguetter",
"mackor",
"drive-in",
"baguette",
"mat",
"gatukök",
"restaurang",
"takeaway",
"bukfylla",
"junk-food",
"bargett",
"fralla",
"frallor",
"grill"
],
"amenity/ferry_terminal":[
"Färjeterminal / Färjehållplats / Färjestation"
],
"amenity/fire_station":[
"brandstång",
"brandbil",
"räddningstjänsten",
"Brandstation",
"brandtorn"
],
"amenity/food_court":[
"mat",
"gatukök",
"mattorg",
"restaurangtorg",
"snabbmat",
"food court",
"restaurang",
"Restaurangtorg"
],
"amenity/fountain":[
"springbrunn",
"Fontän",
"vattenkonst"
],
"amenity/fuel":[
"bensin",
"diesel",
"LNG",
"Bensinstation",
"bränsle",
"propan",
"tapp",
"tankstation",
"CNG",
"mack",
"biodiesel"
],
"amenity/grave_yard":[
"Gravplats",
"urnlund",
"griftegård",
"kyrkogård",
"begravningsplats",
"Kyrkogård",
"minneslund"
],
"amenity/grit_bin":[
"sand",
"Sandlåda",
"salt",
"halkbekämpning",
"Sandkista",
"sandkista",
"sandbehållare",
"halka"
],
"amenity/hospital":[
"sanatorium",
"sjukhus",
"läkare",
"Sjukhusområde",
"klinik",
"sjukvård",
"institution",
"lasarett",
"läkarmottagning",
"sjukstuga",
"vårdhem",
"kirurgi",
"sjuk"
],
"amenity/hunting_stand":[
"jakt",
"skjuta",
"viltjakt",
"Jakttorn",
"utkik",
"älgtorn",
"utkikstorn",
"vilt",
"Skjutstege"
],
"amenity/ice_cream":[
"glasskiosk",
"yogurt",
"glass",
"Glassaffär",
"mjukglass",
"sorbet",
"sherbet",
"frozen",
"kulglass",
"gelato"
],
"amenity/internet_cafe":[
"Internetcafé",
"internetkafé",
"internetcaffe",
"internetcafe",
"cybercafé",
"Internetkafé"
],
"amenity/kindergarten":[
"kindergarten",
"Förskola",
"lekplats",
"Förskoleområde",
"dagis",
"lekskola",
"daghem",
"lekis"
],
"amenity/language_school":[
"språk",
"språkkurs",
"Språkskola",
"språkutbildning",
"esl"
],
"amenity/library":[
"läsesal",
"bokrum",
"Bibliotek",
"boksamling",
"bibbla",
"böcker",
"bokskatt",
"bok"
],
"amenity/love_hotel":[
"Kärlekshotell",
"hotell",
"sexhotell",
"korttidshotell"
],
"amenity/marketplace":[
"Marknadsplats",
"salutorg",
"marknad",
"torg",
"Saluhall"
],
"amenity/monastery":[
"helgedom",
"allah",
"församling",
"tempelområde",
"kyrka",
"katedral",
"religiös anläggning",
"kor",
"vallfärdsort",
"andaktsrum",
"gudshus",
"tillbedjan",
"moské",
"begravningskapell",
"andligt område",
"moske",
"fristad",
"kloster",
"dopkapell",
"kapell",
"gudstjänstslokal",
"tro",
"mission",
"bönehus",
"gud",
"dyrkan",
"guds hus",
"kristendom",
"missionshus",
"sanktuarium",
"andaktssal",
"dom",
"kyrkogård",
"böneplats",
"basilika",
"tempel",
"kyrkobyggnad",
"religiös",
"religiöst område",
"Klosterområde",
"bönhus",
"sidokapell",
"kranskapell",
"predikan",
"vallfärgsplats",
"betel",
"kristen",
"kyrkbyggnad",
"synagoga",
"mässkapell",
"religion",
"annexkyrka",
"gravkapell",
"kyrkorum",
"andaktslokal",
"gudstjänstlokal",
"gudstjänst",
"kyrksal",
"korkapell",
"tabernakel"
],
"amenity/motorcycle_parking":[
"motorcykelställ",
"parkeringsplats",
"ställplats",
"motorcykel",
"parkering motorcykel",
"parkeringsplats motorcykel",
"Motorcykelparkering",
"parkering"
],
"amenity/music_school":[
"musikskola",
"musikinstrument",
"sångskola",
"kultur",
"kör",
"instrument",
"musik",
"kulturskola",
"instrumentskola",
"sång",
"Musikskola"
],
"amenity/nightclub":[
"diskotek",
"dansställe",
"klubb",
"bar",
"nöjeslokal",
"Nattklubb",
"disco",
"disko*",
"dans",
"dansklubb"
],
"amenity/nursing_home":[
"Vårdhem"
],
"amenity/parking":[
"parkeringsplats",
"bil",
"p-plats",
"bilparkering",
"Parkering",
"parkeringsområde",
"Parkeringsplats"
],
"amenity/parking/multi-storey":[
"parkeringsbyggnad",
"flervånig",
"bil",
"Flervånig bilparkering",
"flervånig parkeringsgarage",
"parkeringshus",
"garage",
"bilparkering",
"parkeringsgarage",
"inomhusparkering",
"parkering",
"parkeringsramp",
"parkeringsdäck",
"garagebyggnad",
"Flervånigt parkeringsgarage"
],
"amenity/parking_entrance":[
"utfart",
"garage",
"parkeringshus",
"infart",
"In- och utfart parkeringsgarage"
],
"amenity/parking_space":[
"handikapsparkering",
"handikapsficka",
"Parkeringsruta",
"parkeringsyta",
"Enskild parkeringsplats",
"parkeringsficka"
],
"amenity/pharmacy":[
"Läkemedel",
"drog*",
"medicin",
"Läkemedel*",
"droghandel",
"apotek",
"läkemedelsaffär",
"farmaceut",
"recept"
],
"amenity/place_of_worship":[
"helgedom",
"allah",
"församling",
"tempelområde",
"kyrka",
"katedral",
"religiös anläggning",
"kor",
"vallfärdsort",
"andaktsrum",
"gudshus",
"tillbedjan",
"moské",
"begravningskapell",
"andligt område",
"moske",
"fristad",
"kloster",
"dopkapell",
"kapell",
"gudstjänstslokal",
"tro",
"mission",
"bönehus",
"gud",
"dyrkan",
"guds hus",
"kristendom",
"missionshus",
"sanktuarium",
"andaktssal",
"dom",
"kyrkogård",
"böneplats",
"basilika",
"tempel",
"kyrkobyggnad",
"religiös",
"religiöst område",
"Plats för tillbedjan",
"bönhus",
"sidokapell",
"kranskapell",
"socken",
"predikan",
"vallfärgsplats",
"betel",
"kristen",
"kyrkbyggnad",
"synagoga",
"mässkapell",
"religion",
"slottskapell",
"annexkyrka",
"gravkapell",
"kyrkorum",
"andaktslokal",
"gudstjänstlokal",
"gudstjänst",
"kyrksal",
"korkapell",
"pastorat",
"tabernakel"
],
"amenity/place_of_worship/buddhist":[
"pagoda",
"Buddhisttempel",
"Buddhism",
"Buddha",
"kloster",
"meditation",
"zendo",
"chörten",
"stupa",
"tempel",
"dojo",
"vihara"
],
"amenity/place_of_worship/christian":[
"helgedom",
"församling",
"tempelområde",
"kyrka",
"katedral",
"religiös anläggning",
"kor",
"vallfärdsort",
"andaktsrum",
"gudshus",
"tillbedjan",
"begravningskapell",
"andligt område",
"fristad",
"Kyrka",
"kloster",
"dopkapell",
"kapell",
"gudstjänstslokal",
"tro",
"mission",
"bönehus",
"gud",
"dyrkan",
"guds hus",
"kristendom",
"missionshus",
"sanktuarium",
"andaktssal",
"dom",
"kyrkogård",
"böneplats",
"basilika",
"tempel",
"kyrkobyggnad",
"religiös",
"religiöst område",
"bönhus",
"sidokapell",
"kranskapell",
"socken",
"predikan",
"vallfärgsplats",
"betel",
"kristen",
"kyrkbyggnad",
"mässkapell",
"religion",
"slottskapell",
"annexkyrka",
"gravkapell",
"kyrkorum",
"andaktslokal",
"gudstjänstlokal",
"gudstjänst",
"kyrksal",
"korkapell",
"pastorat",
"tabernakel"
],
"amenity/place_of_worship/hindu":[
"hinduism",
"helgedom",
"hindu",
"Hindutempel",
"garbhagriha",
"Sanatana Dharma",
"puja",
"arcana",
"tempel"
],
"amenity/place_of_worship/jewish":[
"helgedom",
"dom",
"predikan",
"katedral",
"Synagoga",
"böneplats",
"tempel",
"religion",
"Jude",
"tro",
"bönehus",
"gudshus",
"gudstjänstlokal",
"Judendom",
"tillbedjan",
"missionshus"
],
"amenity/place_of_worship/muslim":[
"helgedom",
"muslim",
"predikan",
"böneplats",
"religion",
"kyrkobyggnad",
"tro",
"bönehus",
"gudshus",
"gudstjänstlokal",
"tillbedjan",
"moské",
"minaret",
"Moské"
],
"amenity/place_of_worship/shinto":[
"kami",
"helgedom",
"torii",
"Jinja",
"shintohelgedom",
"shrine",
"tempel",
"yashiro",
"jingū",
"Shinto shrine",
"miya",
"Shinto",
"Jinja (Shintoistisk helgedom)",
"shintoism"
],
"amenity/place_of_worship/sikh":[
"helgedom",
"Sikh-tempel",
"Sikh",
"Sikhtempel",
"Sikhism",
"Gurudwara",
"Sikhiskt tempel",
"tempel"
],
"amenity/place_of_worship/taoist":[
"helgedom",
"Taoistiskt tempel",
"Taoism",
"tao",
"daoism",
"tempel"
],
"amenity/planetarium":[
"museum",
"observatorium",
"astronomi",
"Planetarium"
],
"amenity/police":[
"polisman",
"pass",
"poliskonstapel",
"Polis",
"snut",
"polismyndighet",
"kriminalare",
"ordningsmakt",
"polisväsende",
"lag",
"konstapel",
"polismakt",
"polisstation"
],
"amenity/post_box":[
"Postlåda",
"brevinkast",
"post",
"Brevlåda",
"postlåda",
"brev"
],
"amenity/post_office":[
"Postkontor",
"post",
"kort",
"postverk",
"posten",
"frimärke",
"paket",
"försändelser",
"postgång",
"postväsende",
"brev"
],
"amenity/prison":[
"häkte",
"fångvårdsanstalt",
"polisarrest",
"Fängelseområde",
"fängelse",
"arrest",
"anstalt",
"fängelseförvar",
"fånganstalt",
"finka"
],
"amenity/pub":[
"bar",
"ölservering",
"nattklubb",
"öl",
"sprit",
"alkohol",
"ölstuga",
"drinkar",
"Pub",
"krog"
],
"amenity/public_bath":[
"badinrättning",
"het källa",
"badhus",
"simbassäng",
"bad",
"bassängbad",
"bassäng",
"badplats",
"strandbad",
"onsen",
"strand",
"Publikt bad",
"fotbad",
"badställe"
],
"amenity/public_bookcase":[
"begagnade böcker",
"Offentlig bokhylla",
"publik bokhylla",
"låneböcker",
"bokdelning",
"bibliotek",
"bokbyte"
],
"amenity/ranger_station":[
"informationscenter",
"infocenter",
"besökscenter",
"friluftsområde",
"Friluftsanläggningen",
"park",
"friluftsliv"
],
"amenity/recycling":[
"Återvinning"
],
"amenity/recycling_centre":[
"skräp",
"återvinningsstation",
"flaskor",
"dumpa",
"Återvinningscentral",
"glas",
"sopstation",
"skrot",
"återbruk",
"burkar",
"återvinning",
"sopor"
],
"amenity/recycling_container":[
"skräp",
"container",
"metall",
"återvinningscontainer",
"återvinningsstation",
"flaskor",
"glas",
"återbruk",
"Återvinningscontainer ",
"sopstation",
"skrot",
"burkar",
"återvinning",
"sopor"
],
"amenity/register_office":[
"Registreringsbyrå"
],
"amenity/restaurant":[
"café. matsal",
"lunch",
"servering",
"grillbar",
"värdshus",
"kafé",
"brasserie",
"cafeteria",
"krog",
"bodega",
"rotisseri",
"matservering",
"bar",
"matställe",
"pizzeria",
"Restaurang",
"restauration",
"pub",
"näringsställe",
"sylta",
"kaffe"
],
"amenity/restaurant/american":[
"lunch",
"servering",
"grillbar",
"värdshus",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"matställe",
"näringsställe",
"kaffe",
"café. matsal",
"USA",
"kafé",
"amerikansk mat",
"bodega",
"rotisseri",
"pizzeria",
"Restaurang",
"restauration",
"pub",
"amerikansk restaurang",
"sylta",
"Amerikansk restaurang"
],
"amenity/restaurant/asian":[
"café. matsal",
"asiatisk restaurang",
"lunch",
"servering",
"grillbar",
"värdshus",
"kafé",
"brasserie",
"cafeteria",
"krog",
"bodega",
"rotisseri",
"matservering",
"bar",
"matställe",
"Asiatisk restaurang",
"pizzeria",
"asiatisk mat",
"Restaurang",
"restauration",
"pub",
"näringsställe",
"sylta",
"kaffe"
],
"amenity/restaurant/chinese":[
"lunch",
"servering",
"grillbar",
"värdshus",
"kinesisk",
"kinesisk restaurang",
"brasserie",
"cafeteria",
"kinamat",
"krog",
"matservering",
"bar",
"Kina",
"Kinesisk restaurang",
"matställe",
"näringsställe",
"kaffe",
"café. matsal",
"kafé",
"bodega",
"rotisseri",
"pizzeria",
"Restaurang",
"restauration",
"pub",
"sylta"
],
"amenity/restaurant/french":[
"fransk restaurang",
"lunch",
"servering",
"Frankrike",
"grillbar",
"värdshus",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"matställe",
"Fransk restaurang",
"näringsställe",
"kaffe",
"café. matsal",
"kafé",
"bodega",
"rotisseri",
"pizzeria",
"Restaurang",
"restauration",
"pub",
"fransk mat",
"sylta"
],
"amenity/restaurant/german":[
"lunch",
"servering",
"grillbar",
"värdshus",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"matställe",
"tysk mat",
"näringsställe",
"kaffe",
"tysk restaurang",
"café. matsal",
"Tyskland",
"kafé",
"Tysk restaurang",
"bodega",
"rotisseri",
"pizzeria",
"Restaurang",
"restauration",
"pub",
"sylta"
],
"amenity/restaurant/greek":[
"Grekisk restaurang",
"lunch",
"servering",
"grillbar",
"värdshus",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"matställe",
"grekisk restaurang",
"näringsställe",
"kaffe",
"café. matsal",
"grekisk mat",
"kafé",
"bodega",
"rotisseri",
"Grekland",
"pizzeria",
"Restaurang",
"restauration",
"pub",
"sylta"
],
"amenity/restaurant/indian":[
"lunch",
"servering",
"grillbar",
"värdshus",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"matställe",
"indisk restaurang",
"näringsställe",
"kaffe",
"indisk mat",
"café. matsal",
"kafé",
"bodega",
"rotisseri",
"pizzeria",
"Indisk restaurang",
"Restaurang",
"restauration",
"pub",
"Indien",
"sylta"
],
"amenity/restaurant/italian":[
"lunch",
"servering",
"grillbar",
"värdshus",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"matställe",
"Italiensk restaurang",
"näringsställe",
"kaffe",
"café. matsal",
"kafé",
"bodega",
"rotisseri",
"italiensk mat",
"pizzeria",
"Restaurang",
"restauration",
"pub",
"sylta",
"Italien",
"italiensk restaurang"
],
"amenity/restaurant/japanese":[
"lunch",
"servering",
"Japansk restaurang",
"grillbar",
"värdshus",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"matställe",
"näringsställe",
"kaffe",
"café. matsal",
"japansk restaurang",
"Japan",
"kafé",
"bodega",
"rotisseri",
"pizzeria",
"japansk mat",
"Restaurang",
"restauration",
"pub",
"sylta"
],
"amenity/restaurant/mexican":[
"lunch",
"servering",
"grillbar",
"värdshus",
"mexikansk restaurang",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"matställe",
"näringsställe",
"kaffe",
"café. matsal",
"Mexiko",
"Mexikansk restaurang",
"kafé",
"bodega",
"rotisseri",
"pizzeria",
"mexikansk mat",
"Restaurang",
"restauration",
"pub",
"sylta"
],
"amenity/restaurant/noodle":[
"lunch",
"servering",
"grillbar",
"värdshus",
"risnudlar",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"matställe",
"nudlar",
"ris",
"näringsställe",
"kaffe",
"café. matsal",
"Nudelrestaurang",
"kafé",
"nudelrestaurang",
"bodega",
"rotisseri",
"pizzeria",
"Restaurang",
"restauration",
"pub",
"sylta"
],
"amenity/restaurant/pizza":[
"lunch",
"servering",
"grillbar",
"värdshus",
"brasserie",
"cafeteria",
"krog",
"pan-pizza",
"matservering",
"bar",
"matställe",
"pizza",
"panpizza",
"näringsställe",
"kaffe",
"café. matsal",
"pan pizza",
"pizzarestaurang",
"kafé",
"bodega",
"rotisseri",
"pizzeria",
"Restaurang",
"restauration",
"pub",
"Pizzarestaurang",
"sylta"
],
"amenity/restaurant/seafood":[
"hummer",
"lunch",
"kräftdjur",
"servering",
"grillbar",
"värdshus",
"blötdjur",
"Fisk- och skaldjursrestaurang",
"brasserie",
"cafeteria",
"krog",
"krabba",
"fiskerestaurang",
"matservering",
"bar",
"matställe",
"bläckfisk",
"näringsställe",
"kaffe",
"café. matsal",
"seafood",
"kafé",
"bodega",
"skaldjur",
"rotisseri",
"räkor",
"skaldjursrestaurang",
"fisk",
"ostron",
"krabbor",
"pizzeria",
"Restaurang",
"restauration",
"pub",
"sylta",
"musslor"
],
"amenity/restaurant/steakhouse":[
"lunch",
"servering",
"grillbar",
"värdshus",
"steakhouse",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"matställe",
"steak house",
"näringsställe",
"kaffe",
"kött",
"café. matsal",
"Stekhus",
"biff",
"kafé",
"bodega",
"rotisseri",
"pizzeria",
"Restaurang",
"restauration",
"pub",
"slakthus",
"sylta",
"stekhus"
],
"amenity/restaurant/sushi":[
"lunch",
"servering",
"grillbar",
"värdshus",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"matställe",
"asiatisk mat",
"sushi",
"näringsställe",
"kaffe",
"café. matsal",
"asiatisk restaurang",
"kafé",
"bodega",
"rotisseri",
"Sushi-restaurang",
"pizzeria",
"Restaurang",
"restauration",
"pub",
"sylta"
],
"amenity/restaurant/thai":[
"lunch",
"servering",
"grillbar",
"värdshus",
"Thai-restaurang",
"brasserie",
"cafeteria",
"Thailand",
"krog",
"matservering",
"bar",
"matställe",
"asiatisk mat",
"thaimat",
"näringsställe",
"kaffe",
"café. matsal",
"asiatisk restaurang",
"thai",
"kafé",
"bodega",
"rotisseri",
"pizzeria",
"Restaurang",
"restauration",
"pub",
"sylta"
],
"amenity/restaurant/turkish":[
"lunch",
"servering",
"grillbar",
"värdshus",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"matställe",
"Turkiet",
"näringsställe",
"kaffe",
"café. matsal",
"Turkisk restaurang",
"kafé",
"bodega",
"rotisseri",
"turkisk mat",
"turkisk",
"pizzeria",
"Restaurang",
"restauration",
"pub",
"sylta"
],
"amenity/restaurant/vietnamese":[
"lunch",
"servering",
"grillbar",
"värdshus",
"brasserie",
"cafeteria",
"krog",
"matservering",
"bar",
"Vietnam",
"matställe",
"asiatisk mat",
"Vietnamesisk restaurang",
"Vietnamesisk mat",
"näringsställe",
"kaffe",
"café. matsal",
"asiatisk restaurang",
"kafé",
"bodega",
"rotisseri",
"pizzeria",
"Restaurang",
"restauration",
"pub",
"sylta"
],
"amenity/sanitary_dump_station":[
"tömningsplats",
"gråvatten",
"toalettömning",
"Campingtoalett",
"sanitet",
"campingplats",
"torrtoalett",
"Latrintömning"
],
"amenity/school":[
"Campus",
"högskoleområde",
"gymnasium",
"grundskola",
"Skolområde",
"universitet",
"Skolgård",
"högskola",
"högstadium",
"mellanstadium",
"universitetsområde",
"skolområde",
"lågstadium"
],
"amenity/scrapyard":[
"Bilskrot"
],
"amenity/shelter":[
"väntkur",
"grotta",
"hydda",
"Skydd",
"vindskydd",
"Väderskydd",
"koja",
"väderskydd",
"tak över huvudet",
"picknick",
"lusthus"
],
"amenity/shelter/gazebo":[
"trädgårdspaviljong",
"fåfänga",
"paviljong",
"Lusthus",
"kolonistuga"
],
"amenity/shelter/lean_to":[
"gapskjul",
"Vindskydd",
"skärmskydd"
],
"amenity/shelter/picnic_shelter":[
"Picknicktak",
"Picknickplats",
"rastplats",
"paviljong",
"pavilion",
"utflykt",
"Picknick"
],
"amenity/shelter/public_transport":[
"busskur",
"busshållplats",
"väntplats",
"skydd",
"väderskydd",
"spårvagnshållplats",
"Väderskydd för kollektivtrafik"
],
"amenity/shower":[
"duschbad",
"Dusch",
"duschrum",
"badrum",
"duschkabin",
"duschutrymme"
],
"amenity/smoking_area":[
"rökruta",
"cigarett",
"Rökområde",
"rökning tillåten",
"rökrum",
"röka",
"rökning",
"rökområde"
],
"amenity/social_facility":[
"uteliggare",
"social",
"välgörenhetsorganisationer",
"social hjälp",
"socialen",
"välgörenhet",
"hjälparbete",
"Social inrättning"
],
"amenity/social_facility/food_bank":[
"matbank",
"Matbank",
"välgörenhetsorganisation",
"matutdelning",
"matpaket"
],
"amenity/social_facility/group_home":[
"grupphem",
"välgörenhetsorganisationer",
"gammal",
"välgörenhet",
"hjälparbete",
"ålderdomshem",
"Gruppboende",
"kollektiv"
],
"amenity/social_facility/homeless_shelter":[
"Härbärge",
"hemlös",
"sovsal",
"bostadslös"
],
"amenity/social_facility/nursing_home":[
"pensionärshem",
"servicehus",
"hem för gamla",
"Seniorboende",
"servicehem",
"äldreboende",
"HVB-hem",
"seniorboende",
"senior",
"pensionär",
"assistansboende",
"Vårdhem",
"ålderdomshem",
"hem för vård och boende"
],
"amenity/studio":[
"utsändningslokal",
"TV",
"filminspelning",
"inspelningslokal",
"television",
"TV-studio",
"inspelning",
"filmstudio",
"Studio",
"radiostudio",
"radio"
],
"amenity/swimming_pool":[
"Simbassäng"
],
"amenity/taxi":[
"taxificka",
"taxistation",
"taxi",
"Taxihållplats"
],
"amenity/telephone":[
"telefonautomat",
"telefonkiosk",
"telefonkur",
"telefonhytt",
"Telefon"
],
"amenity/theatre":[
"skådebana",
"drama",
"Teater",
"teaterföreställning",
"föreställning",
"skådespel",
"skådeplats",
"scen",
"musikal",
"pjäs",
"teater"
],
"amenity/theatre/type/amphi":[
"utomhus",
"utomhusteater",
"läktare",
"scen",
"Amfiteater",
"teater",
"utescen"
],
"amenity/toilets":[
"avträde",
"latrin",
"Toalett",
"hemlighus",
"skithus",
"badrum",
"toa",
"Toaletter",
"utedass",
"bekvämlighetsinrättning",
"wc",
"Baja-Maja",
"klo",
"vattentoalett",
"dass",
"torrklosett",
"klosett",
"vattenklosett",
"bajamaja",
"mugg"
],
"amenity/townhall":[
"ämbetsverk",
"folkets hus",
"Stadshus",
"fullmäktige",
"riksdag",
"domstolsbyggnad",
"parlament",
"samlingslokal",
"myndighet",
"representation",
"samlingsplats",
"stad",
"Kommunhus",
"kommunalhus",
"by",
"kommun",
"kommunstyrelse",
"förvaltning"
],
"amenity/university":[
"college",
"universitetsbyggnad",
"högskola",
"högskoleområde",
"Universitet",
"universitetsområde",
"akademi",
"Universitetsområde",
"lärosäte"
],
"amenity/vehicle_inspection":[
"Bilbesiktning",
"Fordonsbesiktning",
"bilprovningen",
"fordonsinspektion",
"Bilprovning",
"besiktning",
"bilinspektion"
],
"amenity/vending_machine":[
"biljett",
"tuggummiautomater",
"läsk",
"Varuautomat",
"biljettautomat",
"läskautomat",
"varumaskin",
"biljetter",
"godisautomat",
"mellanmål"
],
"amenity/vending_machine/cigarettes":[
"cigaretter",
"snusautomat",
"tobaksautomat",
"Cigarettautomat"
],
"amenity/vending_machine/coffee":[
"the",
"te",
"Varuautomat",
"Espresso",
"expresso",
"Kaffeautomat",
"varumaskin",
"kaffe"
],
"amenity/vending_machine/condoms":[
"kondomomat",
"Kondomautomat",
"kondomer"
],
"amenity/vending_machine/drinks":[
"kaffeautomat",
"drickautomat",
"läsk",
"dryck",
"dryckesautomat",
"Dryckesautomat ",
"läskautomat",
"kaffemaskin",
"juice",
"kaffe",
"dryckautomat"
],
"amenity/vending_machine/electronics":[
"kabel",
"laddare",
"kablar",
"varumaskin",
"laddkabel",
"laddkablar",
"mobiltelefon",
"pekplatta",
"telefon",
"surfplatta",
"varuautomat",
"Varumaskin för elektronik",
"elektronik",
"öronsnäckor",
"hörlurar"
],
"amenity/vending_machine/elongated_coin":[
"mynt",
"Penny Press",
"minnesmyntmaskin",
"elongated penny",
"myntpressmaskin",
"ECM",
"coin maskin",
"minne",
"minnesmynt",
"souvenirmynt",
"elongated coin-maskin",
"Elongated coin-maskin (myntpressmaskin)",
"elongated coin",
"souvenir"
],
"amenity/vending_machine/excrement_bags":[
"hundpåsar",
"hund",
"bajs",
"hundskit",
"Bajspåsar",
"hundbajs",
"avföringspåse",
"djur",
"skitpåse",
"hundbajspåsar"
],
"amenity/vending_machine/feminine_hygiene":[
"Varumaskin för mensskydd",
"kvinnor",
"binda",
"tampong",
"kvinna",
"bindor",
"menstruation",
"kondom",
"mens",
"mensskydd"
],
"amenity/vending_machine/food":[
"mat",
"matvarumaskin",
"matautomat",
"Matvaruautomat",
"Varuautomat",
"varumaskin",
"mellanmål"
],
"amenity/vending_machine/fuel":[
"Bränslepump",
"diesel",
"ing",
"tanka",
"bensinstation",
"propan",
"tankomat",
"tankstation",
"mack",
"bensin",
"etanol",
"bränsle",
"tapp",
"pump",
"cng",
"biodiesel"
],
"amenity/vending_machine/ice_cream":[
"glass",
"Glassautomat",
"Varuautomat",
"isglass",
"varumaskin"
],
"amenity/vending_machine/news_papers":[
"Tidningsautomat"
],
"amenity/vending_machine/newspapers":[
"Tidningsautomat",
"tidning",
"tidningsdistribution",
"tidningar",
"tidningsutlämning",
"tidningslåda"
],
"amenity/vending_machine/parcel_pickup":[
"amazon",
"webbshop",
"paketutlämning",
"leverans",
"internetbutik",
"InPosts",
"paketautomat",
"paketleverans",
"paket",
"utlämning",
"Paketautomat (utlämning)"
],
"amenity/vending_machine/parcel_pickup_dropoff":[
"amazon",
"packetinlämning",
"webbshop",
"paketutlämning",
"leverans",
"internetbutik",
"InPosts",
"paketautomat",
"paketleverans",
"paket",
"utlämning",
"Paketautomat (ut- och inlämning)"
],
"amenity/vending_machine/parking_tickets":[
"parkeringsur",
"biljett",
"parkeringsavgift",
"parkometer",
"Parkeringsautomat",
"parkering"
],
"amenity/vending_machine/public_transport_tickets":[
"tågbiljett",
"tågbiljetter",
"transport",
"tunnelbana",
"färja",
"båt",
"Biljettautomat för kollektivtrafik",
"bussbiljetter",
"biljett",
"tåg",
"bussbiljett",
"spårvagn",
"Biljettautomat",
"buss"
],
"amenity/vending_machine/stamps":[
"porto",
"frankering",
"post",
"Varuautomat",
"Frimärksautomat",
"frankeringsautomat",
"varumaskin",
"frimärke",
"vykort",
"brev"
],
"amenity/vending_machine/sweets":[
"tuggummi",
"tuggummiautomater",
"chips",
"godis",
"Godisautomat",
"godisautomat",
"mellanmål"
],
"amenity/veterinary":[
"djurdoktor",
"djurläkare",
"djurklinik",
"Veterinär ",
"djursjukhus",
"Veterinär"
],
"amenity/waste/dog_excrement":[
"hund",
"sopkärl",
"hundbajspåse",
"bajs",
"Sopkärl för hundbajspåsar",
"hundskit",
"hundbajs",
"bajspåsar",
"skitpåse",
"hundbajspåsar",
"soptunna"
],
"amenity/waste_basket":[
"skräpkorg",
"skräp",
"Soptunna",
"Soptunna (liten)",
"sopkärl",
"papperskorg",
"papperskärl",
"avfallskorg",
"sopor"
],
"amenity/waste_disposal":[
"Soptunna",
"industrisopor",
"sopkärl",
"avfall",
"avfallskärl",
"avfallstunna",
"hushållssopor",
"avfallskontainer",
"Soptunna (hushålls- eller industrisopor)",
"sopor"
],
"amenity/waste_transfer_station":[
"skräp",
"dumpa",
"skrot",
"återvinning",
"Avfallscentral"
],
"amenity/water_point":[
"Dricksvatten",
"vattenpåfyllning",
"Dricksvatten för campingfordon"
],
"amenity/watering_place":[
"dricksvatten",
"utfodring",
"dricksvatten för djur",
"djurutfodring",
"Dricksvatten för djur",
"vattenhåll",
"djur",
"vattenkar"
],
"area":[
"fällt",
"areal",
"område",
"utrymme",
"Yta",
"plan",
"mark"
],
"area/highway":[
"vägplan",
"Vägbeläggning",
"Vägyta",
"torg",
"köryta",
"promenatyta"
],
"attraction/amusement_ride":[
"karusell",
"Åkattraktion",
"nöjespark",
"temapark",
"tivoli",
"nöjeskarusell"
],
"attraction/animal":[
"akvarium",
"lejon",
"björn",
"Djur",
"apa",
"temapark",
"djurpark",
"fiskar",
"zoo",
"tiger",
"zoologisk trädgård"
],
"attraction/big_wheel":[
"åkattraktion",
"karusell",
"nöjespark",
"temapark",
"stort hjul",
"tivoli",
"Pariserhjul",
"nöjeskarusell"
],
"attraction/bumper_car":[
"åkattraktion",
"Radiobilar",
"nöjespark",
"temapark",
"radiobil",
"tivoli"
],
"attraction/bungee_jumping":[
"Bungyjump",
"bungee jump",
"nöjespark",
"temapark",
"hopplattform",
"tivoli"
],
"attraction/carousel":[
"åkattraktion",
"nöjespark",
"temapark",
"Karusell",
"Karusell (roterande)",
"tivoli",
"nöjeskarusell"
],
"attraction/dark_ride":[
"åkattraktion",
"karusell",
"nöjespark",
"temapark",
"tivoli",
"spöktåg",
"Mörk åktur",
"nöjeskarusell"
],
"attraction/drop_tower":[
"åkattraktion",
"karusell",
"nöjespark",
"temapark",
"tivoli",
"Fritt fall",
"nöjeskarusell"
],
"attraction/maze":[
"Trojeborg",
"slingergång",
"Trädgårdslabyrint",
"Labyrint",
"Trojaborg",
"irrgång"
],
"attraction/pirate_ship":[
"karusell",
"roterande båt",
"vikingaskepp",
"Åkattraktion",
"nöjespark",
"temapark",
"gunga",
"tivoli",
"Båtgunga",
"piratskepp",
"gungande båt",
"nöjeskarusell"
],
"attraction/river_rafting":[
"karusell",
"Åkattraktion",
"nöjespark",
"temapark",
"forsbana",
"fors",
"tivoli",
"Forsränning",
"Vattenbana",
"nöjeskarusell"
],
"attraction/roller_coaster":[
"åkattraktion",
"berg- och dalbana",
"bergochdalbana",
"dalbana",
"Berg- och dalbana",
"nöjespark",
"temapark",
"berg-och-dalbana",
"berg-och-dal-bana",
"bergodalbana",
"tivoli"
],
"attraction/summer_toboggan":[
"kälke",
"Sommarrodel",
"rodel",
"Sommerrodelbahn",
"mountain coaster",
"Alpine slide"
],
"attraction/train":[
"stadståg",
"sightseeing",
"vägtåg",
"sightseeingtåg",
"Turisttåg (ej på räls)",
"turisttåg",
"Tschu-Tschu",
"Tuff tuff-tåg"
],
"attraction/water_slide":[
"vattenrutschkana",
"Vattenrutschbana",
"rutschkana",
"vattenrutschbana"
],
"barrier":[
"bom",
"räcke",
"avspärrning",
"stopp",
"Barriär",
"skydd",
"hinder",
"blockering",
"mur",
"barriär",
"vall",
"spärr"
],
"barrier/block":[
"trafikbarriärer",
"sugga",
"Block",
"Trafikhinder",
"betongsugga",
"avspärrare"
],
"barrier/bollard":[
"Pollare",
"stolpe",
"Stolpe"
],
"barrier/border_control":[
"passkontroll",
"pass",
"tull",
"Gränskontroll",
"säkerhetskontroll",
"gräns"
],
"barrier/cattle_grid":[
"Färist",
"galler",
"rist"
],
"barrier/city_wall":[
"skans",
"vallar",
"Stadsmur",
"befästningsverk",
"fort",
"barrikad",
"mur",
"ringmur"
],
"barrier/cycle_barrier":[
"Cykelbarriär",
"Cykelbarriär ",
"hinder",
"barriär"
],
"barrier/ditch":[
"ränna",
"Dike",
"vallgrav"
],
"barrier/entrance":[
"Entré"
],
"barrier/fence":[
"gärdsgård",
"inhägnad",
"stängsel",
"Staket"
],
"barrier/gate":[
"Grind"
],
"barrier/hedge":[
"Häck",
"buskar"
],
"barrier/kerb":[
"trottoarkant",
"kantsten",
"Trottoarkant",
"kant"
],
"barrier/kerb/lowered":[
"trottoarkant",
"kantsten",
"Nedsänkt trottoarkant",
"sluttande",
"nedsänkt trottoar",
"barnvagnsramp",
"kantstensramp",
"trottoarsramp",
"rullstolsramp",
"kantstensskärning",
"kant",
"nedsänkt kant"
],
"barrier/kissing_gate":[
"Grind vid betesmark",
"Kryssgrind"
],
"barrier/lift_gate":[
"Bom",
"avspärrning",
"lyftbom",
"spärr"
],
"barrier/retaining_wall":[
"Stödmur",
"nivåskillnad"
],
"barrier/stile":[
"Övergång",
"trappa"
],
"barrier/toll_booth":[
"vägavgift",
"importavgift",
"tullmyndighet",
"gränstull",
"tullvisitation",
"tullkontroll",
"Tullstation",
"tullhus",
"införselavgift",
"skatt"
],
"barrier/wall":[
"befästning",
"vägg",
"hinder",
"murverk",
"Mur",
"skyddsvärn",
"barriär"
],
"boundary/administrative":[
"Gräns",
"gränslinje",
"Administrativ gräns",
"administrativ gräns"
],
"bridge/support":[
"pylon",
"stödpelarna",
"anfang",
"bropelare",
"landfäste",
"akvedukt",
"Brostöd",
"snedkabelbro",
"stöd",
"viadukt",
"förankring",
"hängbro",
"bro"
],
"bridge/support/pier":[
"akvedukt",
"stöd",
"viadukt",
"vägport",
"överfart",
"stödpelare",
"pelare",
"balkbro",
"bro",
"Stödpelare"
],
"building":[
"anläggning",
"fastighet",
"kåk",
"bygge",
"konstruktion",
"hus",
"Byggnad",
"byggnadsverk"
],
"building/barn":[
"lagård",
"loge",
"ladugård",
"Lada",
"magasin",
"skjul",
"skulle"
],
"building/boathouse":[
"Båthus",
"sjöbod",
"strandbod"
],
"building/bungalow":[
"fristående hus",
"stuga",
"sommarstuga",
"Bungalow",
"semesterhus",
"villa"
],
"building/bunker":[
"Bunker"
],
"building/cabin":[
"kåk",
"Stuga",
"sommarstuga",
"hus",
"koja",
"fritidshus",
"landställe",
"torp"
],
"building/carport":[
"Carport",
"garage",
"bilparkering",
"biltak",
"övertäckt parkering",
"parkering"
],
"building/cathedral":[
"helgedom",
"dom",
"stiftskyrka",
"Katedral",
"kyrka",
"religiös anläggning",
"kyrkogård",
"basilika",
"kyrkobyggnad",
"Huvudkyrka",
"religiös",
"religiöst område",
"vallfärdsort",
"gudshus",
"biskopskyrka",
"tillbedjan",
"andligt område",
"fristad",
"kloster",
"predikan",
"vallfärgsplats",
"kristen",
"kyrkbyggnad",
"religion",
"tro",
"kyrkorum",
"gud",
"biskop",
"dyrkan",
"guds hus",
"gudstjänst",
"kyrksal",
"domkyrka",
"kristendom"
],
"building/chapel":[
"helgedom",
"andaktssal",
"tempelområde",
"kyrka",
"religiös anläggning",
"kyrkogård",
"böneplats",
"kor",
"tempel",
"kyrkobyggnad",
"religiös",
"religiöst område",
"bönhus",
"sidokapell",
"andaktsrum",
"gudshus",
"tillbedjan",
"begravningskapell",
"fristad",
"socken",
"predikan",
"dopkapell",
"kristen",
"Kapell",
"kyrkbyggnad",
"mässkapell",
"religion",
"tro",
"slottskapell",
"gravkapell",
"annexkyrka",
"kyrkorum",
"mission",
"bönehus",
"andaktslokal",
"gudstjänstlokal",
"gud",
"Kranskapell",
"dyrkan",
"guds hus",
"gudstjänst",
"kyrksal",
"korkapell",
"kristendom",
"missionshus",
"sanktuarium"
],
"building/church":[
"helgedom",
"församling",
"tempelområde",
"katedral",
"religiös anläggning",
"kor",
"vallfärdsort",
"gudshus",
"andaktsrum",
"tillbedjan",
"begravningskapell",
"andligt område",
"fristad",
"Kyrka",
"kloster",
"dopkapell",
"kapell",
"gudstjänstslokal",
"tro",
"mission",
"bönehus",
"gud",
"dyrkan",
"guds hus",
"Kyrkobyggnad",
"kristendom",
"missionshus",
"sanktuarium",
"andaktssal",
"dom",
"kyrkogård",
"böneplats",
"basilika",
"tempel",
"kyrkobyggnad",
"religiös",
"religiöst område",
"bönhus",
"sidokapell",
"kranskapell",
"socken",
"predikan",
"vallfärgsplats",
"betel",
"kristen",
"kyrkbyggnad",
"mässkapell",
"religion",
"slottskapell",
"annexkyrka",
"gravkapell",
"kyrkorum",
"andaktslokal",
"gudstjänst",
"kyrksal",
"korkapell",
"pastorat",
"tabernakel"
],
"building/civic":[
"kommunal",
"stadshus",
"kommunhus",
"Civil",
"publik",
"Kommunal byggnad",
"medborgarhus"
],
"building/college":[
"Gymnasie",
"gymnasium",
"gymnasiebyggnad",
"Collegebyggnad",
"universitet"
],
"building/commercial":[
"Kommersiell byggnad",
"kommersiellt",
"Kontorsbyggnad",
"affärsbyggnad",
"handelsbyggnad"
],
"building/construction":[
"bygge",
"byggarbete",
"byggnadsplats",
"byggarbetsplats",
"byggnation",
"Byggnad under uppförande",
"Byggnad under konstruktion"
],
"building/detached":[
"enfamiljshus",
"fristående hus",
"Villa",
"hus",
"friliggande villa",
"Fristående hus",
"friliggande hus",
"envåningshus",
"fristående villa",
"egnahem",
"kåk",
"enbostadshus",
"småhus"
],
"building/dormitory":[
"sovsal",
"Elevhem",
"korridorboende",
"internatskola",
"internat",
"kollektiv",
"Korridorboende",
"studentkorridor"
],
"building/entrance":[
"Entré/utgång"
],
"building/farm":[
"lantbruk",
"gård",
"Mangårdsbyggnad",
"bostadshus",
"hus",
"Mangårdsbyggnad (bostadshus på gård)",
"bostad"
],
"building/farm_auxiliary":[
"lantbruk",
"ekonomibyggnader",
"gård",
"ladugård",
"gårdshus",
"stall",
"Gårdsbyggnader",
"lantbruksbyggnader"
],
"building/garage":[
"kallgarage",
"Garage",
"bilskjul",
"garage",
"parkeringshus",
"varmgarage",
"bilstall",
"carport"
],
"building/garages":[
"kallgarage",
"bilgarage",
"Garage",
"bilförvaring",
"bilskjul",
"parkeringshus",
"uppställningsplats",
"varmgarage",
"bilstall",
"skydd för bilar",
"carport"
],
"building/grandstand":[
"åskådarplats",
"åskådare",
"Huvudläktare",
"sittplats",
"läktare",
"publik",
"sport"
],
"building/greenhouse":[
"vinterträdgård",
"Växthus",
"driveri",
"blomsterhus",
"orangeri",
"odlingshus",
"växthus",
"drivhus",
"växtodling"
],
"building/hospital":[
"sjukvårdsinrättning",
"klinik",
"lasarett",
"sjukhem",
"sjukstuga",
"vårdhem",
"sjukhus",
"Sjukhusbyggnad",
"hospital",
"vårdanstalt"
],
"building/hotel":[
"",
"motell",
"hotell",
"Hotellbyggnad",
"vandrarhem",
"värdshus",
"härbärge",
"pensionat",
"gästhem"
],
"building/house":[
"enfamiljshus",
"kåk",
"Villa",
"bostadshus",
"enbostadshus",
"hus",
"småhus",
"Enfamiljshus",
"parhus",
"egnahem",
"radhus"
],
"building/hut":[
"barack",
"hydda",
"stuga",
"skydd",
"Koja",
"kyffe"
],
"building/industrial":[
"lager",
"Industribyggnad",
"industri",
"fabrik"
],
"building/kindergarten":[
"dagishus",
"förskolehus",
"kindergarten",
"förskolebyggnad",
"Förskola",
"barnomsorg",
"dagis",
"lekskola",
"dagisbyggnad",
"daghem",
"lekis",
"Förskolebyggnad"
],
"building/mosque":[
"Moskébyggnad",
"islam",
"muslim",
"muhammedansk helgedom",
"muhammedanism",
"moské",
"minaret"
],
"building/pavilion":[
"Klubbhus",
"Sport",
"omklädningsrum",
"paviljong",
"klubbhus",
"idrott",
"idrottsklubb"
],
"building/public":[
"allmän byggnad",
"offentlig byggnad",
"Publik byggnad"
],
"building/residential":[
"Hyreshus",
"Boningshus",
"Bostadshus",
"Flerfamiljshus"
],
"building/retail":[
"Affärsbyggnad",
"detaljhandel",
"butik",
"försäljningsställe",
"varuhus",
"kiosk",
"affärshus",
"affärer"
],
"building/roof":[
"överbyggnad",
"valv",
"övertäckning",
"regnskydd",
"Tak"
],
"building/ruins":[
"husrest",
"fornlämning",
"raserad",
"förfallen",
"ödehus",
"huslämning",
"ruin",
"Ruinbyggnad"
],
"building/school":[
"gymnasium",
"skolhus",
"undervisning",
"grundskola",
"utbildning",
"skola",
"undervisningsanstalt",
"högstadium",
"folkhögskola",
"mellanstadium",
"komvux",
"Skolbyggnad",
"läroanstalt",
"läroverk",
"skolväsen",
"lärosäte",
"lågstadium"
],
"building/semidetached_house":[
"fristående hus",
"Villa",
"radhusområde",
"hus",
"friliggande hus",
"småhus",
"parhus",
"Delvist Fristående hus",
"radhus",
"parhusområde"
],
"building/service":[
"teknikhus",
"transformator",
"nätstation",
"Teknikhus",
"teknik",
"transformatorhus",
"fördelningsstation",
"mäthus",
"pumphus",
"mätstation",
"pump",
"mätning"
],
"building/shed":[
"uthus",
"förråd",
"visthusbod",
"visthus",
"Skjul",
"förvaring",
"verkstad",
"förvaringsskjul",
"barack",
"hobbyhus",
"bod",
"friggebod",
"hobbyrum"
],
"building/stable":[
"stallbyggnad",
"hästar",
"ridhusanläggning",
"ridhus",
"Stall",
"häst"
],
"building/stadium":[
"arenabyggnad",
"stadion",
"byggnad",
"Stadionbyggnad",
"friidrottsstadion",
"stadium",
"Stadion",
"arena"
],
"building/static_caravan":[
"husvagn",
"campingvagn",
"Villavagn"
],
"building/temple":[
"fristad",
"helgedom",
"tempelområde",
"religiös anläggning",
"böneplats",
"tempel",
"religion",
"tro",
"religiös",
"religiöst område",
"Tempelbyggnad",
"mission",
"bönehus",
"bönhus",
"andaktsrum",
"gudshus",
"gud",
"dyrkan",
"guds hus",
"tillbedjan"
],
"building/terrace":[
"Terrasshus"
],
"building/train_station":[
"Järnvägsstation"
],
"building/transportation":[
"Byggnad för kollektivtrafik",
"linbaneterminal",
"Färjeterminal",
"linbana",
"linjetrafik",
"terminal",
"transport",
"färja",
"båt",
"kollektivtrafikbyggnad",
"kollektivtrafik",
"Perrong",
"bussterminal",
"båtterminal",
"spårvagnsterminal",
"metro",
"transit",
"station",
"buss"
],
"building/university":[
"högskola",
"Universitetsbyggnad",
"högskolebyggnad",
"universitet"
],
"building/warehouse":[
"lager",
"lada",
"upplag",
"depå",
"packhus",
"Lagerhus",
"magasin"
],
"camp_site/camp_pitch":[
"tält",
"camping",
"husvagn",
"Tältplats/husvagnsplats",
"Campingplats",
"husvagnsplats",
"Tältplats"
],
"circular":[
"Trafikcirkel"
],
"club":[
"klubblokal",
"klubb",
"föreningslokal",
"förening",
"Klubb",
"sammanslutning",
"socialt",
"sällskap"
],
"craft":[
"hantverkare",
"Hantverk",
"skrå",
"slöjd"
],
"craft/basket_maker":[
"korgflätning",
"korgtillverkning",
"Korgtillverkare",
"korg",
"Korgslöjd"
],
"craft/beekeeper":[
"honung",
"bi",
"honungstillverkning",
"Biodlare",
"biodling"
],
"craft/blacksmith":[
"konsthantverk",
"smide",
"smidesverkstad",
"smida",
"Smed"
],
"craft/boatbuilder":[
"båtbyggeri",
"varv",
"båtbyggare",
"Båtbyggare"
],
"craft/bookbinder":[
"bokbinderi",
"bokbindning",
"bindning",
"Bokbindare",
"böcker",
"bokreparatör",
"bok"
],
"craft/brewery":[
"ölframställning",
"öl",
"Bryggeri",
"öltillverkning"
],
"craft/carpenter":[
"timmerman",
"byggnadssnickare",
"träarbetare",
"grovsnickare",
"Snickare"
],
"craft/carpet_layer":[
"matta",
"mattläggning",
"golv",
"golvläggare",
"Mattläggare"
],
"craft/caterer":[
"matleverantör",
"matleverans",
"catering",
"Catering",
"cateringfirma"
],
"craft/chimney_sweeper":[
"Sotare",
"skorstensfejare",
"rökgång",
"sotarmurre",
"skorsten"
],
"craft/clockmaker":[
"Urmakare (väggur)",
"klockmakare",
"Urmakare"
],
"craft/confectionery":[
"konfekt",
"sötsaker",
"godisfabrik",
"choklad",
"Godistillverkare",
"godis",
"godsaker",
"konfektyrer",
"karameller",
"pastiller"
],
"craft/distillery":[
"sprittillverkning",
"mezcal",
"bourbon",
"alkohol",
"sprit",
"gin",
"hembränning",
"rom",
"tequila",
"whisky",
"vodka",
"alkoholtillverkning",
"spritdryck",
"Destilleri",
"spritdestillering",
"brandy",
"alkoholdestillering",
"scotch"
],
"craft/dressmaker":[
"Sömmerska",
"Dressmaker",
"sy",
"kvinnokläder",
"klädtillverkning",
"skräddare",
"Klädsömmare",
"sömnad",
"klänning",
"kläder"
],
"craft/electrician":[
"systembyggare",
"kabeldragning",
"montör",
"el",
"elkraft",
"elmontör",
"elreparatör",
"starkströmsmontör",
"Elektriker"
],
"craft/electronics_repair":[
"tv-service",
"tv-reparatör",
"datorreparation",
"reparation",
"skärmbyte",
"datorservice",
"telefonreparatör",
"elektronikreparation",
"reparatör",
"elektronik",
"Elektronikreparatör",
"vitvaror",
"tvättmaskinsreparatör"
],
"craft/gardener":[
"landskapsarkitekt",
"Trädgårdsmästare",
"trädgård",
"handelsträdgård"
],
"craft/glaziery":[
"Glasmästare",
"glasblåsare",
"glas",
"fönster",
"solskydd",
"glaskonst",
"målat glas"
],
"craft/handicraft":[
"snickeri",
"hantverk",
"konsthantverk",
"textil",
"Hantverkare",
"vävstuga",
"Hantverk",
"handarbete",
"sömnad",
"slöjd",
"snideri",
"hemslöjd",
"vävning"
],
"craft/hvac":[
"inomhusklimat",
"energiförsörjning",
"ventilation",
"sanitet",
"avlopp",
"kyla",
"VVS",
"värme",
"air condition",
"rörmokare",
"övervakningssystem",
"styrsystem",
"gas",
"vattenförsörjning",
"uppvärmning",
"luftkonditionering",
"tryckluft",
"vatten",
"sprinkler",
"installationsteknik"
],
"craft/insulator":[
"Isolering",
"ljudisolering",
"isolerare",
"värmeisolering",
"isolationsmaterial"
],
"craft/jeweler":[
"Smycken"
],
"craft/key_cutter":[
"nyckelringar",
"Nyckeltillverkning",
"hänglås",
"nyckel",
"nycklar",
"nyckelkopiering",
"nyckelring"
],
"craft/locksmith":[
"Låssmed"
],
"craft/metal_construction":[
"Metallarbete",
"metallarbetare",
"metallindustri",
"kallbearbetning",
"svets",
"svetsare",
"svetsning"
],
"craft/optician":[
"Optiker"
],
"craft/painter":[
"Målare",
"färg",
"måleriarbetare",
"penslar",
"tapetsering",
"måleri",
"tapetserare",
"lackering",
"målarmästare",
"tapeter"
],
"craft/photographer":[
"Fotograf",
"bild",
"fotografering",
"porträttfotografering",
"bildkonst",
"porträtt",
"kamera"
],
"craft/photographic_laboratory":[
"mörkrum",
"Fotoframkallning",
"kanvas",
"framkallning",
"fotoframkallning",
"foto",
"Filmframkallning",
"film",
"utskrift"
],
"craft/plasterer":[
"puts",
"Putsare",
"cement",
"gips",
"väggputs"
],
"craft/plumber":[
"rörmontör",
"rörläggare",
"Rörmokare",
"dränering",
"vatten",
"avlopp",
"rör"
],
"craft/pottery":[
"lergods",
"Krukmakeri",
"krukgods",
"keramik",
"Krukmakare",
"porslin",
"stengods",
"glasering",
"lerkärl",
"drejare",
"drejning",
"lera",
"krukmakeri",
"keramiker"
],
"craft/rigger":[
"tackling",
"rigg",
"segelbåt",
"segelfartyg",
"mast",
"segel",
"Riggare",
"tågvirke"
],
"craft/roofer":[
"Takläggare, takläggning, tak, takpannor, yttertak, Taktegel, tegel",
"Takläggare"
],
"craft/saddler":[
"läder",
"säte",
"Sadelmakare",
"sadelmakeri",
"sadel"
],
"craft/sailmaker":[
"Segelmakare",
"segelsömnad",
"segel",
"segelmakeri"
],
"craft/sawmill":[
"Sågverk",
"trä",
"virke",
"brädor",
"bräda",
"timmer",
"plank"
],
"craft/scaffolder":[
"ställning",
"Ställningsbyggare",
"byggnadsställning"
],
"craft/sculptor":[
"skulptör",
"bildhuggare",
"skulpturer",
"Skulptör",
"bildsnidare",
"skulptur",
"staty"
],
"craft/shoemaker":[
"Skomakare",
"skor"
],
"craft/stonemason":[
"Stenhuggare",
"stenbrott"
],
"craft/tailor":[
"Skräddare"
],
"craft/tiler":[
"golvläggare",
"Plattläggare"
],
"craft/tinsmith":[
"plåtslagare",
"Tennsmed ",
"tenn",
"förtennare",
"Tennsmed",
"Tunnplåtslagare"
],
"craft/upholsterer":[
"Möbelstoppare",
"stoppning",
"tapetserare",
"möbler"
],
"craft/watchmaker":[
"Urmakare (små klockor)",
"Urmakare",
"armbandsur",
"fickur",
"klockreparatör"
],
"craft/window_construction":[
"fönsterinstallatör",
"Fönstertillverkare",
"dörr",
"dörrleverantör",
"dörrar",
"glas",
"dörrmontör",
"dörrinstallatör",
"fönster",
"fönsterleverantör",
"fönstermontör",
"dörrtillverkare"
],
"craft/winery":[
"Vinfabrik",
"vinframställnig",
"vineri",
"vinproduktion",
"Vinframställning",
"vin"
],
"embankment":[
"Vägbank"
],
"emergency/ambulance_station":[
"Ambulansstation",
"räddning",
"räddningstjänst",
"ambulans"
],
"emergency/defibrillator":[
"hjärtstartare",
"Defibrillator",
"hjärthjälp"
],
"emergency/designated":[
"Åtkomst för utryckningsfordon – Avsedd för"
],
"emergency/destination":[
"Åtkomst för utryckningsfordon – Destination"
],
"emergency/fire_alarm":[
"brandtelefon",
"Nödtelefon"
],
"emergency/fire_extinguisher":[
"skumsläckare",
"pulversläckare",
"vattensläckare",
"vattenpost",
"eldsläckare",
"koldioxidsläckare",
"brandsläckning",
"Brandpost",
"Brandsläckare",
"brandslang",
"handbrandsläckare",
"kolsyresläckare",
"brand"
],
"emergency/fire_hydrant":[
"brandsläckning",
"Brandpost",
"vattenpost",
"brandslang"
],
"emergency/first_aid_kit":[
"brännsår",
"sårvård",
"plåster",
"sår",
"Första hjälpen",
"första hjälpen låda",
"första hjälpen kit",
"förbandslåda",
"förband",
"bandage"
],
"emergency/life_ring":[
"livräddningsboj",
"frälsarkrans",
"Livboj",
"livräddning",
"livboj"
],
"emergency/lifeguard":[
"Badvakt",
"CPR",
"strandvakt",
"livräddare",
"badvakt",
"räddning",
"Lifeguard"
],
"emergency/no":[
"Åtkomst för utryckningsfordon – Nej"
],
"emergency/official":[
"Åtkomst för utryckningsfordon – Officiellt"
],
"emergency/phone":[
"nödnummer",
"Nödtelefon",
"alarmtelefon",
"larmtelefon",
"alarmeringscentral"
],
"emergency/private":[
"Åtkomst för utryckningsfordon – Privat"
],
"emergency/siren":[
"larm",
"Viktigt Meddelande till Allmänheten",
"beredskapslarm",
"mistlur",
"starktonssiren",
"varning",
"flyglarm",
"Siren",
"Tyfon",
"Hesa Fredrik",
"VMA"
],
"emergency/water_tank":[
"vattensamling",
"kris",
"reservoar",
"räddning",
"vattentorn",
"nödtank",
"brandsläckningstank",
"lagringstank",
"brandsläckning",
"cistern",
"Vattentank för brandsläckning",
"tank",
"brand",
"nöd",
"vatten",
"vattentank"
],
"emergency/yes":[
"Åtkomst för utryckningsfordon – Ja"
],
"entrance":[
"entré",
"huvudentré",
"dörr",
"utgång",
"Ingång",
"In-/Utgång"
],
"ford":[
"vad",
"Vadställe",
"övergångsställe"
],
"golf/bunker":[
"golf",
"sandhål",
"sandfälla",
"hinder",
"Bunker",
"sandgrop"
],
"golf/fairway":[
"golf",
"Fairway"
],
"golf/green":[
"puttinggreen",
"golf",
"green",
"hål",
"Green"
],
"golf/hole":[
"golf",
"Golfhål",
"hål"
],
"golf/lateral_water_hazard_area":[
"golf",
"vattenhinder",
"out of bounds",
"Oändligt vattenhinder/sidovattenhinder",
"Oändligt vattenhinder",
"sidovattenhinder"
],
"golf/lateral_water_hazard_line":[
"golf",
"vattenhinder",
"out of bounds",
"Oändligt vattenhinder/sidovattenhinder",
"Oändligt vattenhinder",
"sidovattenhinder"
],
"golf/rough":[
"Ruff",
"ruffen",
"ruff",
"gräs"
],
"golf/tee":[
"golf",
"utslagsplats",
"Tee"
],
"golf/water_hazard_area":[
"golf",
"Vattenhinde"
],
"golf/water_hazard_line":[
"golf",
"Vattenhinde"
],
"healthcare":[
"klinik",
"institution",
"välmående",
"Hälsovård",
"doktor",
"sjukdom",
"kirurgi",
"sjuk",
"läkare",
"hälsa",
"mottagning"
],
"healthcare/alternative":[
"naturopati",
"reiki",
"tuina",
"hydroterapi",
"herbalism",
"antroposofisk",
"hypnos",
"unani",
"ayurveda",
"Alternativmedicin",
"aromaterapi",
"osteopati",
"shiatsu",
"tillämpad kinesiologi",
"örtmedicin",
"homeopati",
"reflexologi",
"traditionell",
"alternativ medicin",
"akupunktur"
],
"healthcare/alternative/chiropractic":[
"ryggen",
"ryggsmärta",
"ryggrad",
"ryggbesvär",
"smärta",
"Kiropraktor",
"Kiropraktik",
"Kiropraktik (rygg)",
"Kotknackare"
],
"healthcare/audiologist":[
"hörapparat",
"Audionom",
"Audionomist",
"Audionomi (hörsel)",
"Audionomi",
"öra",
"örat",
"hörsel",
"ljud"
],
"healthcare/birthing_center":[
"BB",
"graviditet",
"barnafödsel",
"Förlossning",
"bäbis",
"barn",
"Förlossningsavdelning",
"baby",
"förlossning",
"Barnbördshus ",
"bebis"
],
"healthcare/blood_donation":[
"blodgivning",
"blodcentral",
"plasmaferes",
"donera blod",
"blodtransfusion",
"bloddonation",
"ge blod",
"stamcellsdonation",
"Blodgivarcentral",
"blodgivare",
"aferes",
"Plateletpheresis",
"blodbank"
],
"healthcare/hospice":[
"Hospis",
"döende",
"död",
"Palliativ vård",
"terminalvård",
"Hospis (palliativ vård)"
],
"healthcare/laboratory":[
"Medicinskt laboratorium",
"diagnos",
"kemi",
"blodkontroll",
"diagnosering",
"lab",
"immunologi",
"Laboratoriemedicin",
"patologi",
"laboratorium",
"analys",
"medicinskt laboratorium",
"provtagning",
"genetik",
"farmakologi",
"analysrådgivning",
"mikrobiologi",
"blodanalys",
"medicinskt lab",
"transfusionsmedicin"
],
"healthcare/midwife":[
"mödrahälsovård",
"ungdomsmottagning",
"Gynekologi",
"gynekolog",
"jordemo",
"ackuschörska",
"Preventivmedel",
"Barnmorska",
"mödravårdscentra"
],
"healthcare/occupational_therapist":[
"ergonomi",
"terapeut",
"Arbetsterapi",
"rehabilitering",
"hjälpmedel",
"terapi"
],
"healthcare/optometrist":[
"korrektionsglas",
"ögon",
"glasögon",
"Optometri (ögon)",
"Optometrier",
"Optometri",
"linser",
"syn",
"synhjälpmedel",
"synfel",
"ögonlaser"
],
"healthcare/physiotherapist":[
"Fysioterapi (sjukgymnastik)",
"terapeut",
"sjukgymnastik",
"Fysioterapi",
"fysisk",
"Fysioterapeut",
"terapi"
],
"healthcare/podiatrist":[
"Podiatri (fötter)",
"fötter",
"fothälsa",
"fotkirurgi",
"Podiatri",
"naglar",
"podiatriker",
"fot"
],
"healthcare/psychotherapist":[
"Psykoterapi",
"terapeut",
"rådgivare",
"psykolog",
"Psykoterapeut",
"sinne",
"ångest",
"kuratorer",
"självmord",
"terapi",
"psykologisk behandling",
"mental hälsa",
"depression"
],
"healthcare/rehabilitation":[
"Rehabilitering",
"Rehab",
"terapeut",
"terapi"
],
"healthcare/speech_therapist":[
"röst",
"språk",
"terapeut",
"Logoped (röst/tal)",
"dysfagi",
"Logoped",
"språkstörning",
"röststörning",
"tal",
"terapi",
"talstörning"
],
"highway":[
"Väg"
],
"highway/bridleway":[
"rida",
"ryttare",
"ridstig",
"Ridväg",
"ridning",
"häst"
],
"highway/bus_guideway":[
"guidad buss",
"Spårbuss",
"buss"
],
"highway/bus_stop":[
"Busshållplats / Bussplattform"
],
"highway/corridor":[
"inomhus",
"inomhuskorridor",
"korridor",
"gång",
"gångpassage",
"förbindelsegång",
"Korridor inomhus"
],
"highway/crossing/marked":[
"Vägövergång",
"vägpassage",
"gångpassage",
"Markerad gångpassage",
"övergångsställe",
"gångvägspassage",
"Övergångsställe för gående",
"markerat övergångsställe"
],
"highway/crossing/marked-raised":[
"Markerat övergångsställe (upphöjt)",
"Vägövergång",
"vägpassage",
"puckel",
"Övergångsställe för gående",
"markerat övergångsställe",
"gångpassage",
"Markerad gångpassage",
"Markerad gångpassage (upphöjt)",
"fartpuckel",
"fartgupp",
"farthinder",
"övergångsställe",
"gångvägspassage",
"gupp"
],
"highway/crossing/unmarked":[
"Omarkerad gångpassage",
"Omarkerad övergång",
"Vägövergång",
"vägpassage",
"gångpassage",
"övergångsställe",
"gångvägspassage",
"Övergångsställe för gående",
"omarkerat övergångsställe"
],
"highway/crossing/unmarked-raised":[
"Vägövergång",
"vägpassage",
"omarkerat övergångsställe (upphöjt)",
"puckel",
"Övergångsställe för gående",
"omarkerat övergångsställe",
"Omarkerad övergång (upphöjt)",
"Omarkerad övergång",
"gångpassage",
"fartpuckel",
"fartgupp",
"farthinder",
"övergångsställe",
"gångvägspassage",
"gupp"
],
"highway/crossing/zebra":[
"Markerat övergångsställe"
],
"highway/crossing/zebra-raised":[
"Markerat övergångsställe (upphöjt)"
],
"highway/cycleway":[
"cykelled",
"gång- och cykelväg",
"cykelväg",
"gc-väg",
"Cykelväg",
"cykel"
],
"highway/elevator":[
"Hiss"
],
"highway/footway":[
"gång- och cykelväg",
"vandring",
"gångväg",
"gc-väg",
"vandra",
"stig",
"Gångväg",
"löparbana",
"motionsspår",
"promenad"
],
"highway/footway/conveying":[
"gångrullband",
"transportband för människor",
"Rullande trottoar",
"transportband",
"rullband",
"rullande gåband",
"rullande trottoar",
"rullramp",
"transportband för personer",
"rullande gångbana",
"Rullgångbana",
"rulltrottoar"
],
"highway/footway/marked":[
"Markerat övergångsställe",
"Vägövergång",
"vägpassage",
"gångpassage",
"Markerad gångpassage",
"övergångsställe",
"gångvägspassage",
"Övergångsställe för gående",
"markerat övergångsställe"
],
"highway/footway/marked-raised":[
"Markerat övergångsställe (upphöjt)",
"Vägövergång",
"vägpassage",
"puckel",
"Övergångsställe för gående",
"markerat övergångsställe",
"gångpassage",
"Markerad gångpassage",
"Markerad gångpassage (upphöjt)",
"fartpuckel",
"fartgupp",
"farthinder",
"övergångsställe",
"gångvägspassage",
"gupp"
],
"highway/footway/sidewalk":[
"Trottoar",
"gångbana",
"gångväg"
],
"highway/footway/unmarked":[
"Omarkerad gångpassage",
"Omarkerad övergång",
"Vägövergång",
"vägpassage",
"gångpassage",
"övergångsställe",
"gångvägspassage",
"Övergångsställe för gående",
"omarkerat övergångsställe"
],
"highway/footway/unmarked-raised":[
"Vägövergång",
"vägpassage",
"omarkerat övergångsställe (upphöjt)",
"puckel",
"Övergångsställe för gående",
"omarkerat övergångsställe",
"Omarkerad övergång (upphöjt)",
"Omarkerad övergång",
"gångpassage",
"fartpuckel",
"fartgupp",
"farthinder",
"övergångsställe",
"gångvägspassage",
"gupp"
],
"highway/footway/zebra":[
"Markerat övergångsställe"
],
"highway/footway/zebra-raised":[
"Markerat övergångsställe (upphöjt)"
],
"highway/give_way":[
"utfartsregeln",
"lämna företräde",
"väjningspliktsskylt",
"utfart",
"väjningsplikt",
"Väjningsplikt",
"företräde"
],
"highway/living_street":[
"torg",
"Gångfartsområde",
"gårdsgata"
],
"highway/milestone":[
"milstolpe",
"Väghållningsten",
"postament",
"Milsten"
],
"highway/mini_roundabout":[
"Minirondell",
"cirkulationsplats",
"rondell",
"trafikrondell"
],
"highway/motorway":[
"Motorväg",
"snabbled",
"stadsmotorväg"
],
"highway/motorway_junction":[
"motorvägspåfart",
"trafikplats",
"mot",
"avfart",
"Motorvägspåfart / -avfart",
"motorvägsavfart",
"Påfart",
"vägkorsning"
],
"highway/motorway_link":[
"trafikplats",
"motorvägsanslutning",
"avfart",
"Anslutning",
"påfart",
"Anslutning, motorväg"
],
"highway/passing_place":[
"passage",
"Mötesplats",
"passeringsplats",
"möte"
],
"highway/path":[
"vandring",
"gångväg",
"gång",
"vandra",
"vandringsled",
"Stig",
"led",
"spår",
"löparbana",
"motionsspår",
"promenad"
],
"highway/pedestrian_area":[
"plaza",
"gångområde",
"centrum",
"gångväg",
"torg",
"gångfart",
"Gångfartsområde",
"Gågateområde",
"gågata",
"gårdsgata"
],
"highway/pedestrian_line":[
"gångområde",
"affärsgata",
"centrum",
"gångväg",
"gång",
"gående",
"torg",
"shoppinggata",
"promenad",
"plaza",
"gångbana",
"Gågata",
"fotgängare"
],
"highway/primary":[
"primärväg",
"riksväg",
"Primär väg",
"länsväg",
"huvudväg"
],
"highway/primary_link":[
"Anslutning, primär väg",
"primärväg",
"avfart",
"riksväg",
"primär väg",
"Anslutning",
"påfart",
"huvudväg"
],
"highway/raceway":[
"racerbana",
"motorbana",
"gokart",
"rallybana",
"motorracerbana",
"go-kart",
"Motorracerbana",
"tävlingsbana",
"motortävling",
"rally",
"kappkörning"
],
"highway/residential":[
"bostadsområde",
"Bostadsgata",
"gata",
"villaväg",
"villagata"
],
"highway/rest_area":[
"bensinstation",
"Rastplats"
],
"highway/road":[
"främmande",
"ospecificerad",
"Okänd väg",
"okänd väg",
"okänd",
"obekant",
"outforskad"
],
"highway/secondary":[
"sekundärväg",
"länsväg",
"Sekundär väg",
"huvudväg"
],
"highway/secondary_link":[
"sekundär väg",
"Anslutning, sekundär väg",
"avfart",
"sekundärväg",
"länsväg",
"Anslutning",
"påfart",
"huvudväg"
],
"highway/service":[
"Serviceväg",
"bakgård",
"campinggata",
"parkeringsväg",
"Uppfart",
"industriväg"
],
"highway/service/alley":[
"Gränd",
"bigata",
"gränd",
"sidogata",
"bakgata"
],
"highway/service/drive-through":[
"hämtmat",
"McDrive",
"Drive-through",
"Genomkörning"
],
"highway/service/driveway":[
"privat väg",
"garageinfart",
"Uppfart",
"infart",
"villaväg"
],
"highway/service/emergency_access":[
"räddningsväg",
"brandbil",
"nödväg",
"Brandväg",
"polis",
"utrymningsväg",
"brandkår",
"Utryckningsfordon",
"ambulans",
"utryckningsväg",
"Åtkomst för utryckningsfordon"
],
"highway/service/parking_aisle":[
"parkeringsplats",
"Parkeringsväg",
"parkeringsgata"
],
"highway/services":[
"bensinstation",
"snabbmat",
"restaurang",
"Rastplats",
"vägmat",
"Rastplats med försäljning"
],
"highway/speed_camera":[
"fartkontroll",
"hastighetskamera",
"Trafiksäkerhetskamera",
"Fartkamera"
],
"highway/steps":[
"rulltrappa",
"trappor",
"trapp",
"Trappa",
"trappsteg",
"trappnedgång",
"trappuppgång"
],
"highway/steps/conveying":[
"Rulltrappa",
"trappa",
"rörlig trappa"
],
"highway/stop":[
"lämna företräde",
"stopp",
"Stoppskylt"
],
"highway/street_lamp":[
"lyktstolpe",
"Gatlampa ",
"lampa",
"Gatubelysning",
"belysning",
"gatuljus",
"Gatlampa"
],
"highway/tertiary":[
"Tertiär väg",
"sekundära länsväg",
"huvudgata",
"allmän väg",
"länsväg"
],
"highway/tertiary_link":[
"huvudgata",
"Anslutning, tertiär väg",
"avfart",
"länsväg",
"Anslutning",
"påfart",
"tertiär väg"
],
"highway/track":[
"jordbruksväg",
"Jordbruks-/skogsväg",
"åkerväg",
"traktor",
"timmer",
"brandväg",
"jordbruk",
"brandgata",
"virkesväg",
"Bruksväg",
"skogsmaskin",
"åker",
"traktorväg",
"skogsväg",
"timmerväg"
],
"highway/traffic_mirror":[
"utfartspegel",
"spegel",
"hörn",
"konvex",
"Trafikspegel",
"vägspegel",
"säkerhet"
],
"highway/traffic_signals":[
"trafikljus",
"Trafikljus",
"signalljus",
"Trafiksignaler",
"trafiksignal",
"ljus",
"stoppljus"
],
"highway/trunk":[
"riksväg",
"Huvudväg",
"Europaväg",
"motortrafikled"
],
"highway/trunk_link":[
"avfart",
"Europaväg",
"Anslutning, huvudväg",
"Anslutning",
"påfart",
"huvudväg"
],
"highway/turning_circle":[
"Vändplan",
"vändplats",
"Vändplats",
"återvändsgata"
],
"highway/turning_loop":[
"refug",
"Vändslinga (refug)",
"Vändslinga",
"vändlop",
"vändplats"
],
"highway/unclassified":[
"mindre väg",
"Mindre/oklassificerad väg",
"övrig väg",
"Oklassificerad väg",
"industrigata",
"enskild väg",
"skogsväg",
"liten väg",
"industriväg"
],
"historic":[
"Historisk plats",
"historia",
"arv",
"historik"
],
"historic/archaeological_site":[
"historia",
"utgrävning",
"Arkeologisk plats",
"ruin",
"arkeologi",
"historisk plats"
],
"historic/boundary_stone":[
"Gränsmärke",
"Gränssten",
"milsten",
"råmärke",
"gränsröse"
],
"historic/castle":[
"Slott",
"herrsäte",
"fästning",
"borg",
"palats",
"resident"
],
"historic/memorial":[
"Minnesmärke",
"monument",
"minnessten",
"minnestavla"
],
"historic/monument":[
"Monument",
"Minnesmärke",
"monument"
],
"historic/ruins":[
"husras",
"rest",
"ödehus",
"Ruiner",
"lämning",
"Ruin",
"förfallen byggnad"
],
"historic/tomb":[
"Grav",
"gravhög",
"Mausoleum",
"krigsgrav",
"pyramid",
"klippgrav",
"katakomb",
"massgrav",
"Sarkofag",
"krypta",
"gravvalv"
],
"historic/wayside_cross":[
"kors vid väg",
"Kors vid väg",
"Vägkors",
"pilgrim",
"krucifix"
],
"historic/wayside_shrine":[
"helgedom",
"Helgedom längs väg",
"Helgedom vid väg",
"helgedom vid väg",
"pilgrim"
],
"historic/wreck":[
"båt",
"vrak",
"mast",
"skrov",
"Skeppsvrak",
"skepp"
],
"internet_access/wlan":[
"Surfzon",
"wifi",
"wifi hotspot",
"wi-fi",
"hotspot",
"surfzon",
"trådlöst lokalt nät",
"wi-fi hotspot",
"öppet trådlöst nät",
"wlan",
"trådlöst nät",
"uppkopplingszon",
"fritt trådlöst nät"
],
"junction":[
"vägkorsningar",
"trafikplats",
"gatukorsning",
"Korsning",
"vägkors",
"stoppsignal",
"järnvägskorsning",
"trafiksignal",
"stoppskylt",
"korsning",
"cirkulationsplats",
"trafikkorsning",
"övergångsställe",
"rondell"
],
"landuse":[
"Markanvändning",
"användningsområde",
"landanvändning"
],
"landuse/allotments":[
"odlingslott",
"lott",
"koloniträdgård",
"koloniområde",
"Kolonilott",
"Koloniområde",
"täppa"
],
"landuse/aquaculture":[
"Fiskodling",
"alger",
"musselodling",
"pärlodling",
"vattenbruk",
"Akvakultur",
"akvakultur",
"skaldjur",
"Ostronodling",
"vattenväxter",
"räkor",
"fisk",
"utplantering av fisk"
],
"landuse/basin":[
"infiltrering",
"dagvatten",
"bassäng",
"Avrinningsområde",
"avrinning",
"dagvattenbassäng",
"avrinningsområde",
"infiltration"
],
"landuse/brownfield":[
"Brownfield",
"rivningstomt",
"byggtomt",
"rivet",
"förorenat",
"industri",
"Industriområde",
"Övergivet industriområde (Brownfield)",
"övergivet",
"ödetomt"
],
"landuse/cemetery":[
"gravfält",
"grav",
"griftegård",
"Gravfällt",
"begravningsplats",
"Kyrkogård"
],
"landuse/churchyard":[
"religiös",
"religiöst område",
"gravkapell",
"kyrkområde",
"kyrka",
"Kyrkogård (utan gravar)",
"kristen",
"begravningskapell",
"Kyrkogård",
"andligt område",
"kristendom",
"religion"
],
"landuse/commercial":[
"Kommersiell",
"shoppingområde",
"handelsområde",
"handel",
"Kommersiell område",
"kommersiellt",
"butiksområde",
"affärsområde"
],
"landuse/construction":[
"Byggarbetsplats",
"bygge",
"byggarbete",
"byggnadsplats",
"byggnation",
"Byggnad under uppförande",
"Byggnad under konstruktion"
],
"landuse/farm":[
"Åkermark"
],
"landuse/farmland":[
"åkerfält",
"lantbruk",
"gärde",
"inäga",
"odlingsfält",
"Åker",
"åkerlapp",
"åkerjord",
"Åkermark",
"odling",
"fält",
"teg",
"åkermark"
],
"landuse/farmyard":[
"lantbruk",
"gård",
"jordbruk",
"lantegendom",
"Bondgård",
"lantgård"
],
"landuse/forest":[
"dunge",
"skogsvård",
"skogsområde",
"Skog (brukad)",
"Skog",
"skogstrakt",
"träd",
"skogsdunge",
"lund",
"skogsplantering"
],
"landuse/garages":[
"parking",
"kallgarage",
"Garageområde",
"bilskjul",
"garage",
"varmgarage",
"bilstall",
"bilplatser",
"carport"
],
"landuse/grass":[
"refug",
"mittremsa",
"Gräs",
"klippt gräs",
"rondell"
],
"landuse/greenfield":[
"Greenfield",
"framtid",
"Planerad byggnation",
"urbanisering",
"planerad byggnation"
],
"landuse/greenhouse_horticulture":[
"vinterträdgård",
"trädgårdsodling",
"driveri",
"blomsterhus",
"orangeri",
"odlingshus",
"blomma",
"växthus",
"drivhus",
"Växthus för trädgårdsväxter",
"växtodling"
],
"landuse/harbour":[
"båt",
"kaj",
"båtterminal",
"båtplats",
"Hamn",
"marin"
],
"landuse/industrial":[
"fabriksområde",
"Industriområde",
"fabriksdistrikt",
"industricentrum"
],
"landuse/industrial/scrap_yard":[
"metall",
"metallskräp",
"skräp",
"bil",
"fordon",
"bärgning",
"Skrotupplag",
"vrak",
"metallavfall",
"metallåtervinning",
"Bilskrot",
"skrotningsanläggning",
"bildemontering",
"skrot",
"metallskrot",
"skrotupplag"
],
"landuse/industrial/slaughterhouse":[
"Slaktare",
"slakteri",
"ko",
"gris",
"fläsk",
"fjäderfän",
"styckning",
"slaktare",
"styckare",
"kalv",
"slakt",
"chark",
"styckningsanläggning",
"kyckling",
"nötkött",
"slakthus",
"kött"
],
"landuse/landfill":[
"avfallsanläggning",
"tipp",
"Soptipp",
"avskrädeshög",
"återvinningscentral"
],
"landuse/meadow":[
"slåttermark",
"Äng"
],
"landuse/orchard":[
"fruktträd",
"äppelträd",
"fruktträdgård",
"Fruktodling"
],
"landuse/plant_nursery":[
"Plantskola",
"handelsträdgård"
],
"landuse/quarry":[
"stenbrytning",
"täkt",
"sand",
"gruva",
"utgrävning",
"sandtäckt",
"sandtag",
"sten",
"Stenbrott/Sandtag",
"stenbrott"
],
"landuse/railway":[
"spårväg",
"Banområde",
"spårkorridor",
"tåg",
"spårvagn",
"järnvägsområde",
"tågområde",
"tågspår",
"järnväg",
"järnvägskorridor",
"spår"
],
"landuse/recreation_ground":[
"grönområde",
"Rekreationsområde",
"parkanläggning",
"friluftsområde",
"rekreationsområde",
"parkområde",
"trädgård",
"Park"
],
"landuse/religious":[
"helgedom",
"tempelområde",
"kyrka",
"religiös anläggning",
"vallfärgsplats",
"kyrkogård",
"Religiöst område",
"kristen",
"synagoga",
"böneplats",
"religion",
"tempel",
"tro",
"religiös",
"vallfärdsort",
"gud",
"dyrkan",
"tillbedjan",
"moské",
"andligt område",
"kristendom",
"moske"
],
"landuse/residential":[
"lägenhetsområde",
"förort",
"villaområde",
"Bostadsområde",
"miljonområde",
"getto"
],
"landuse/retail":[
"försäljningsområde",
"försäljning",
"shoppingområde",
"handel",
"handelsområde",
"Detaljhandel",
"shoppingcenter",
"affärer",
"affärsområde",
"shopping"
],
"landuse/vineyard":[
"druvor",
"château",
"vineri",
"vinodling",
"vin",
"vindruvor",
"vinframställning",
"vinfält",
"Vingård"
],
"leisure":[
"Nöje",
"fritid",
"tidsfördriv",
"förströelse",
"Fritid",
"ledighet"
],
"leisure/adult_gaming_centre":[
"spelmaskiner",
"spel",
"flipper",
"spelmaskin",
"vuxenspel",
"flipperspel",
"Center för vuxenspel"
],
"leisure/amusement_arcade":[
"spelhall",
"pay-to-play-spel",
"arkadmaskin",
"flipperspel",
"arkadspel",
"Arkadhall",
"spelhus",
"arkadhall",
"arkad",
"spel",
"flipper",
"Spelkonsol",
"körsimulatorer",
"videospel"
],
"leisure/bandstand":[
"bandstand",
"orkester-scen",
"orkesterscen",
"paviljong",
"musikestrad",
"musikscen",
"musikpaviljong",
"estrad",
"musik",
"scen",
"Musikestrad",
"orkester"
],
"leisure/beach_resort":[
"semesteranläggning",
"turist",
"Resort",
"turism",
"turistanläggning",
"badort",
"Strandresort",
"rekreationsort",
"semesterresort",
"hotell",
"strand",
"kurort",
"hotellanläggning"
],
"leisure/bird_hide":[
"fågelskådargömsel",
"utsiktstorn",
"fågeltorn",
"fågelskådningstorn",
"fågelskådare",
"fågelskådartorn",
"Torn/gömsle för fågelskådning",
"Fågelskådning",
"vilttorn"
],
"leisure/bleachers":[
"bänk",
"åskådarplats",
"åskådare",
"sittplats",
"Läktare",
"läktare",
"publik",
"sport"
],
"leisure/bowling_alley":[
"kägelspel",
"Bowlinghall",
"kägelsport",
"Bowlingbana",
"bowlinghall",
"bowling"
],
"leisure/common":[
"fritt tillträde",
"Allmänning",
"öppet område",
"allmän mark"
],
"leisure/dance":[
"rotunda",
"valls",
"foxtrot",
"folkets park",
"bal",
"salsa",
"gammaldans",
"Dansbana",
"swing",
"balsal",
"tango",
"danshus",
"bugg",
"jive"
],
"leisure/dancing_school":[
"danskurs",
"foxtrot",
"vals",
"gamaldans",
"dans",
"salsa",
"swing",
"tiodans",
"tango",
"dansutbildning",
"Dansskola",
"bugg",
"jive"
],
"leisure/dog_park":[
"hund",
"rastgård",
"Hundpark",
"hundgård",
"kennel",
"hundrastgård"
],
"leisure/firepit":[
"Eldstad",
"lägereld",
"eldning",
"brasa",
"campingbrasa",
"lägerplats",
"eldgrop",
"grillplats",
"grill",
"grillning"
],
"leisure/fitness_centre":[
"träning",
"styrketräning",
"gym",
"träningslokal",
"Fitnesscenter",
"Gym / Fitnesscenter",
"konditionsträning",
"motionsinstitut",
"styrketräningslokal"
],
"leisure/fitness_centre/yoga":[
"Yoga studio",
"Yogastudio",
"meditation",
"joga"
],
"leisure/fitness_station":[
"träning",
"motion",
"fitness",
"gym",
"naturgym",
"utegym",
"träningsbana",
"träningsspår",
"Utomhusgym"
],
"leisure/fitness_station/balance_beam":[
"träning",
"motion",
"Balansbom",
"fitness",
"Balansbom (träning)",
"gym",
"naturgym",
"utegym",
"balans",
"Utomhusgym"
],
"leisure/fitness_station/box":[
"hoppövning",
"träning",
"låda",
"motion",
"fitness",
"Träningsplattform/trapsteg",
"hopp",
"plattform",
"utomhusgym",
"gym",
"naturgym",
"utegym"
],
"leisure/fitness_station/horizontal_bar":[
"träning",
"pullup",
"hävräcke",
"motion",
"pull-up",
"utomhusgym",
"naturgym",
"utegym",
"räck",
"bar",
"pull up",
"Räckhäv",
"Räck (träning)",
"fitness",
"gym"
],
"leisure/fitness_station/horizontal_ladder":[
"träna",
"träning",
"pullup",
"motion",
"stege",
"utomhusgym",
"naturgym",
"utegym",
"räck",
"pull up",
"bar",
"Monkey Bars",
"fitness",
"gym",
"Armgång"
],
"leisure/fitness_station/hyperextension":[
"träna",
"Hyperextension",
"träning",
"motion",
"utomhusgym",
"naturgym",
"utegym",
"Ryggsträckare",
"rygg",
"fitness",
"gym",
"Roman Chair",
"rygglyft"
],
"leisure/fitness_station/parallel_bars":[
"träna",
"Barrpress",
"barr",
"träning",
"motion",
"fitness",
"Dips",
"utomhusgym",
"gym",
"naturgym",
"utegym"
],
"leisure/fitness_station/push-up":[
"träna",
"pushup",
"träning",
"Armhävningsstation",
"push up",
"motion",
"fitness",
"utomhusgym",
"armhävning",
"gym",
"naturgym",
"utegym"
],
"leisure/fitness_station/rings":[
"träna",
"träning",
"ringar",
"pullup",
"motion",
"pull-up",
"utomhusgym",
"Ringar",
"naturgym",
"utegym",
"pull up",
"fitness",
"gym"
],
"leisure/fitness_station/sign":[
"träna",
"träning",
"motion",
"fitness",
"utomhusgym",
"gym",
"instruktionsskylt",
"naturgym",
"utegym",
"Träningsinstruktioner",
"skylt"
],
"leisure/fitness_station/sit-up":[
"träna",
"crunch",
"träning",
"motion",
"sit up",
"utomhusgym",
"naturgym",
"utegym",
"sit-up",
"Sit-up-ramp. situp-ramp",
"fitness",
"Situp-ramp",
"gym",
"situp"
],
"leisure/fitness_station/stairs":[
"träna",
"trappor",
"träning",
"hoppövning",
"motion",
"utomhusgym",
"naturgym",
"utegym",
"step up",
"trapp",
"steg",
"fitness",
"hopp",
"trappa",
"plattform",
"Träningstrappa",
"gym"
],
"leisure/garden":[
"odlingslott",
"örtgård",
"Trädgård",
"botanisk trädgård",
"botanik",
"plantering",
"zoologisk trädgård",
"park",
"botanisk"
],
"leisure/golf_course":[
"golf",
"golfcenter",
"Golfbana",
"golfanläggning"
],
"leisure/hackerspace":[
"hackare",
"projekt",
"makerspace",
"hackers",
"lan",
"Hackerspace",
"hackerspace",
"hacklab"
],
"leisure/horse_riding":[
"rida",
"ryttare",
"Ridskola",
"ridhus",
"ridklubb",
"ridning",
"stall",
"hästridning",
"häst",
"häst*"
],
"leisure/ice_rink":[
"Skridskobana ",
"hockey",
"skridsko",
"ishockeybana",
"ishockey",
"isrink",
"Skridskobana",
"ishall",
"isbana",
"skridskohall",
"skridskoåkning",
"konstisbana",
"ishockeyhall",
"curling"
],
"leisure/marina":[
"småbåt",
"båt",
"småbåtshamn",
"yacht",
"segelbåt",
"hamn",
"fritidsbåt",
"gästhamn",
"Marina"
],
"leisure/miniature_golf":[
"miniatyrgolf",
"bangolf",
"äventyrsgolf",
"Minigolf"
],
"leisure/nature_reserve":[
"reservat",
"naturpark",
"naturområde",
"nationalpark",
"Naturreservat",
"naturreservat",
"naturskyddsområde"
],
"leisure/outdoor_seating":[
"ölträdgård",
"al fresco",
"servering",
"beer garden",
"utomhusmatsal",
"restaurang",
"Uteservering",
"café",
"bar",
"utomhus",
"terrass",
"pub",
"glassbar"
],
"leisure/park":[
"grönområde",
"oas",
"nöjesträdgård",
"stadsoas",
"skog",
"gräs",
"skogsmark",
"friluftsområde",
"lund",
"Park",
"plaza",
"gräsmatta",
"lekplats",
"esplanad",
"rekreationsområde",
"plantering",
"trädgård",
"park",
"äng"
],
"leisure/picnic_table":[
"Picknickbord",
"bänk",
"bord",
"matbord",
"utflyktsbord",
"Picknick",
"utebord"
],
"leisure/pitch":[
"stadion",
"fällt",
"idrottsplan",
"sportplats",
"Idrottsplats",
"arena",
"plan",
"idrottsanläggning"
],
"leisure/pitch/american_football":[
"Amerikansk fotbollsplan",
"Amerikansk fotboll",
"football",
"Plan för amerikansk fotboll"
],
"leisure/pitch/badminton":[
"Badmintonbana",
"badminton",
"Badmintonplan",
"fjäderboll"
],
"leisure/pitch/baseball":[
"baseballplan",
"Baseball",
"Baseballplan",
"baseball-plan"
],
"leisure/pitch/basketball":[
"Basketplan",
"basket",
"korgboll"
],
"leisure/pitch/beachvolleyball":[
"beachfotboll",
"beachvolleyplan",
"Beachvolleyboll",
"Beachvolleyhall",
"Beachvolleyplan",
"beachhandboll",
"beachvolley",
"strandvolleyboll",
"volleyboll",
"Beachhall",
"beachplan"
],
"leisure/pitch/boules":[
"pétanque",
"Boule",
"Boule/Bocce-plan",
"lyonnaise",
"Bocce"
],
"leisure/pitch/bowls":[
"Shortmat",
"Bowls",
"Bowlsplan"
],
"leisure/pitch/cricket":[
"kricket",
"Cricket",
"Cricketplan",
"kricketplan"
],
"leisure/pitch/equestrian":[
"rida",
"Ridskola",
"trav",
"ridhus",
"ridklubb",
"Ridområde",
"ridning",
"stall",
"dressyr",
"häst",
"häst*",
"galopp",
"ryttare",
"hästridning",
"hästhoppning"
],
"leisure/pitch/rugby_league":[
"rugby football",
"rugby",
"rugger",
"rugbyplan",
"Rugby League",
"Rugby League-plan"
],
"leisure/pitch/rugby_union":[
"Rugby Union-plan",
"rugby football",
"rugby",
"rugger",
"rugbyplan",
"rugby union"
],
"leisure/pitch/skateboard":[
"Skate Park",
"skateboardramp",
"halfpipe",
"Skateboardpark",
"skateboard"
],
"leisure/pitch/soccer":[
"Fotboll",
"fotbollsplan",
"Fotbollsplan"
],
"leisure/pitch/softball":[
"softball",
"baseboll",
"brännboll",
"Softballplan",
"softballplan",
"boboll"
],
"leisure/pitch/table_tennis":[
"ping pong",
"pingis",
"bordtennis",
"pingpongbord",
"Pingisbord",
"Bordtennisbord",
"pingpong"
],
"leisure/pitch/tennis":[
"Tennisbana",
"tennis",
"tennisplan"
],
"leisure/pitch/volleyball":[
"Volleybollplan",
"beachvolleyboll",
"volleyboll"
],
"leisure/playground":[
"Lekplats",
"lek",
"lekområde",
"klätterställning",
"gunga",
"lekpark"
],
"leisure/resort":[
"semesteranläggning",
"rekreationsort",
"turist",
"semesterresort",
"hotell",
"Resort",
"kurort",
"turism",
"turistanläggning",
"badort",
"hotellanläggning"
],
"leisure/running_track":[
"Kapplöpningsbana",
"löpbana",
"motionsspår",
"Löparbana"
],
"leisure/sauna":[
"kölna",
"badstuga",
"sauna",
"Bastu"
],
"leisure/slipway":[
"Stapelbädd",
"sjösättning",
"båtramp",
"Sjösättningsplats",
"staplar",
"varv",
"docka",
"torrdocka",
"fartygsdocka"
],
"leisure/sports_centre":[
"idrottsplats",
"träning",
"sportanläggning",
"idrottsplan",
"motion",
"träningsanläggning",
"fitnes",
"sportpalats",
"Sportcenter",
"idrottshall",
"Sportcenter / -anläggning",
"gym",
"simhall",
"sporthall",
"idrottsanläggning"
],
"leisure/sports_centre/swimming":[
"badhus",
"simbassäng",
"badhall",
"simning",
"Badanläggning",
"pool",
"tävlingssim",
"simhall",
"bassäng",
"swimmingpool",
"motionssim"
],
"leisure/stadium":[
"Stadium",
"arena"
],
"leisure/swimming_pool":[
"Simbassäng",
"simning",
"pool",
"bassäng",
"swimmingpool",
"simma"
],
"leisure/track":[
"cykeltävling",
"cykellopp",
"kapplöpningsbana",
"travbana",
"Tävlingsbana (Icke motorsport)",
"hundkapplöpning",
"Tävlingsbana",
"löpbana",
"galoppbana",
"hästkapplöpning",
"löpning"
],
"leisure/water_park":[
"vattenland",
"Äventyrsbad / Vattenpark",
"vattenlekpark",
"Äventyrsbad",
"Vattenpark"
],
"line":[
"utsträckning",
"sträcka",
"streck",
"Linje"
],
"man_made":[
"artificiell",
"Människoskapat",
"Människoskapad",
"syntetisk",
"konstgjort",
"onaturlig"
],
"man_made/adit":[
"gruvhål",
"Stollen",
"gruvingång",
"stoll",
"gruva",
"gruvgång",
"horisontell gruvgång",
"Horisontell gruvgång (Stoll)",
"lichtloch",
"dagort",
"sidoort"
],
"man_made/antenna":[
"mobil",
"Antenn",
"mobilmast",
"tv",
"överföring",
"mast",
"sändning",
"radiomast",
"tv-mast",
"kommunikation",
"radio"
],
"man_made/breakwater":[
"fördämning",
"hamnarm",
"Vågbrytare",
"pir",
"vågskydd",
"hamnpir"
],
"man_made/bridge":[
"fällbro",
"akvedukt",
"övergång",
"vridbro",
"viadukt",
"vägport",
"överfart",
"förbindelse",
"spång",
"bro",
"Bro"
],
"man_made/bunker_silo":[
"lager",
"Ensilage",
"spannmålssilo",
"spannmål",
"pressfoder",
"foder",
"fodersilo",
"Plansilo",
"silo",
"djurfoder",
"spannmålslagring"
],
"man_made/chimney":[
"Skorsten",
"rökgång",
"skorsten"
],
"man_made/clearcut":[
"föryngringsavverkning",
"skog",
"hygge",
"trä",
"träd",
"kalhygge",
"Kalhygge",
"timmer",
"avverkning",
"föryngringsyta",
"avskogning",
"Slutavverkning",
"skövlat skogsområde",
"avverkningsområde"
],
"man_made/crane":[
"Kran",
"vinsch",
"travers",
"lyftkran",
"telfer"
],
"man_made/cutline":[
"pipelinegata",
"Snittlinje",
"jaktgata",
"skiljelinje",
"skogssektion",
"Snittlinje i skog",
"pipeline",
"rörgata",
"gränslinje",
"skogsområde",
"brandgata",
"skidspår",
"domän",
"gräns",
"rågång"
],
"man_made/embankment":[
"bank",
"Vägbank",
"Upphöjning",
"barnvall",
"vall"
],
"man_made/flagpole":[
"Flaggstång",
"flagga",
"Flaggstolpe"
],
"man_made/gasometer":[
"Gasklocka",
"gasbehållare",
"gasometer",
"gascistern",
"gas",
"cistern",
"stadsgas",
"naturgas"
],
"man_made/groyne":[
"Hövd, vågbrytare vinkelrätt mot kusten",
"vågbrytare",
"pir",
"erosion",
"hövd",
"erosionsskydd"
],
"man_made/lighthouse":[
"fyrtorn",
"fyrskepp",
"Fyr"
],
"man_made/mast":[
"mobiltelefon torn",
"mobilmast",
"stagas torn",
"överföringsmast",
"antennbärare",
"mobiltelefonmast",
"radiomast",
"sändarmast",
"Mast",
"antenn",
"sändarstation",
"slavsändare",
"kommunikationsmast",
"tv-mast",
"tv-torn",
"kommunikationstorn",
"överföringstorn"
],
"man_made/mast/communication":[
"mobilmast",
"överföringsmast",
"radiomast",
"mast",
"radiotorn",
"sändartorn",
"mobilantenn",
"mobiltelefon",
"radiosändning",
"antenn",
"kommunikationsmast",
"transmissionsmast",
"radioantenn",
"TV-mast",
"Kommunikationsmast",
"TV-torn",
"kommunikationstorn",
"överföringstorn"
],
"man_made/mast/communication/mobile_phone":[
"mobilantenn",
"mobiltelefon",
"mobilmast",
"antenn",
"överföringsmast",
"Mobilmast",
"kommunikationsmast",
"transmissionsmast",
"mast",
"kommunikationstorn",
"överföringstorn"
],
"man_made/mast/communication/radio":[
"radiosändning",
"antenn",
"överföringsmast",
"transmissionsmast",
"radiomast",
"mast",
"radiotorn",
"Radiomast",
"radioantenn",
"sändartorn",
"överföringstorn"
],
"man_made/mast/communication/television":[
"mobilmast",
"TV",
"överföringsmast",
"mast",
"radiomast",
"television",
"sändartorn",
"mobilantenn",
"mobiltelefon",
"antenn",
"kommunikationsmast",
"transmissionsmast",
"radioantenn",
"TV-mast",
"TV-sändning",
"TV-torn",
"kommunikationstorn",
"överföringstorn"
],
"man_made/monitoring_station":[
"Seismolog",
"vattennivå",
"radon",
"väderstation",
"trafik",
"väder",
"luftkvalitet",
"observation",
"övervakningsstation",
"observationsrör",
"Mätstation",
"luftkvalité",
"gps",
"jordbävning",
"trafikmätning",
"seismologi",
"luftmätning",
"mätning",
"ljud"
],
"man_made/observatory":[
"astronomisk",
"astronom",
"Observatorium",
"meteorologisk",
"rymd",
"teleskop"
],
"man_made/petroleum_well":[
"olja",
"oljetorn",
"Oljeborrning",
"Oljeborr",
"oljepump",
"petroleum"
],
"man_made/pier":[
"hamnarm",
"vågbrytare",
"kaj",
"Pir",
"hamnpir"
],
"man_made/pipeline":[
"ledning",
"oljeledning",
"avloppsledning",
"vattenledning",
"rörledning",
"Pipeline"
],
"man_made/pumping_station":[
"vattenpump",
"avloppspump",
"Pumpstation",
"oljepump",
"spillvattenspump",
"pump",
"dräneringspump",
"pumpaggregat"
],
"man_made/silo":[
"lager",
"Ensilage",
"spannmålssilo",
"spannmål",
"pressfoder",
"foder",
"fodersilo",
"silo",
"Silo",
"djurfoder",
"spannmålslagring"
],
"man_made/storage_tank":[
"reservoar",
"Lagringstank",
"vattentorn",
"cistern",
"tank"
],
"man_made/surveillance":[
"övervakningsutrustning",
"bevakningskamera",
"bevakning",
"övervakningskamera",
"Övervakning",
"kamera"
],
"man_made/surveillance/camera":[
"ANPR",
"registreringsskylt",
"webbkamera",
"ALPR",
"vakt",
"övervakning",
"Övervakningskamera",
"video",
"kamera",
"CCTV",
"webcam säkerhetskamera",
"säkerhet"
],
"man_made/survey_point":[
"fixpunkt",
"Trianguleringspunkt",
"triangulering",
"kartritning"
],
"man_made/tower":[
"Torn",
"torn",
"radiotorn"
],
"man_made/tower/communication":[
"mobilmast",
"överföringsmast",
"radiomast",
"mast",
"radiotorn",
"sändartorn",
"mobilantenn",
"mobiltelefon",
"radiosändning",
"antenn",
"kommunikationsmast",
"transmissionsmast",
"radioantenn",
"TV-mast",
"Kommunikationstorn",
"TV-torn",
"kommunikationstorn",
"överföringstorn"
],
"man_made/tower/observation":[
"utsiktstorn",
"observationstorn",
"utsiktspost",
"observationspost",
"Utkikstorn",
"brandtorn"
],
"man_made/wastewater_plant":[
"reningsverk",
"avloppsverk",
"vattenreningsverk",
"Avloppsreningsverk",
"vattenrening",
"avlopp"
],
"man_made/water_tower":[
"vattenreservoar",
"Vattentorn",
"vatten"
],
"man_made/water_well":[
"Brunn",
"källa",
"vattenbrunn",
"grundvatten",
"vattenhål"
],
"man_made/water_works":[
"vattenreningsanläggning",
"vattenreningsverk",
"vatten",
"Vattenverk",
"vattenanläggning"
],
"man_made/watermill":[
"vattenmölla",
"kvarnhjul",
"kvarn",
"Vattenkvarn",
"mölla",
"skovelhjul",
"skvalta",
"skvaltkvarn"
],
"man_made/windmill":[
"Väderkvarn",
"vindmölla",
"kvarn",
"mölla",
"vädemölle",
"vindkraft"
],
"man_made/works":[
"fabriksbyggnad",
"bil",
"bearbetningsanläggning",
"montering",
"monteringsanläggning",
"fabrikstillverkning",
"verkstad",
"Fabrik",
"raffinaderi",
"oljeraffinaderi",
"tillverkning",
"plast",
"industri",
"möbeltillverkning",
"bryggeri",
"bearbetning"
],
"manhole":[
"Brunnslock",
"dagvatten",
"telefoni",
"dagvattenbrunn",
"manhålslucka",
"Rensbrunn",
"Gatubrunn",
"manlucka",
"avlopp",
"telekom",
"Brandpost",
"a-brunn",
"avloppsbrunn",
"brunn",
"manhål"
],
"manhole/drain":[
"dagvattenbrunn",
"smältvatten",
"avloppsvatten",
"regnvatten",
"regn",
"avlopp",
"Dagvattenbrunn",
"Dagvatten",
"dagbrunn",
"spillvatten",
"dränering",
"avrinning",
"avloppsbrunn"
],
"manhole/telecom":[
"telekom",
"Brunnslock",
"tele-brunn",
"gatubrunn",
"Manhålslucka för telekom",
"telefoni",
"manhålslucka",
"manlucka",
"tele",
"brunn",
"manhål"
],
"natural":[
"natur",
"Naturligt",
"naturanvändning",
"naturlig",
"geologi",
"Naturlig",
"skyddsområde"
],
"natural/bare_rock":[
"Kala klippor ",
"klippor",
"berghäll",
"häll",
"kala klippor"
],
"natural/bay":[
"bukt",
"Vik"
],
"natural/beach":[
"strandlinje",
"badstrand",
"flodstrand",
"sandstrand",
"badställe",
"Strand",
"grusstrand",
"badplats"
],
"natural/cave_entrance":[
"grotta",
"bergrum",
"berghåla",
"Grottingång",
"bergsöppning",
"grotthål",
"grottöppning",
"grottsystem"
],
"natural/cliff":[
"klippa",
"klippavsats",
"Klippa",
"terrass",
"stup",
"platå",
"brant",
"bergskam"
],
"natural/coastline":[
"strand",
"kustlinje",
"kustremsa",
"ö",
"kust",
"Kustlinje",
"hav"
],
"natural/fell":[
"fjällandskap",
"trädgräns",
"högfjäll",
"Fjäll"
],
"natural/glacier":[
"landis",
"jökel",
"gletscher",
"ismassa",
"Glaciär"
],
"natural/grassland":[
"Grässlätt",
"gräsfällt",
"äng"
],
"natural/heath":[
"tundra",
"slätt",
"alvar",
"hed",
"kalmark",
"Hed",
"slättmark",
"gräs",
"äng",
"stäpp"
],
"natural/mud":[
"sörja",
"sankmark och sumpmark",
"dy",
"våtmark",
"gegga",
"gyttja",
"Lera",
"lerigt"
],
"natural/peak":[
"kulle",
"höjdpunkt",
"alp",
"berg",
"hjässa",
"klint",
"Bergstopp",
"kalott",
"höjd",
"klätt",
"topp",
"klack"
],
"natural/reef":[
"grund",
"rev",
"Sandbank",
"Rev",
"sandbank",
"undervattensgrund",
"sandrev",
"sand",
"undervattensskär",
"bank",
"korall",
"barriär",
"hav",
"revel",
"korallrev"
],
"natural/ridge":[
"kulle",
"horst",
"kam",
"berg",
"höjd",
"högland",
"bergsområde",
"krön",
"ås",
"bergsrygg",
"Ås"
],
"natural/saddle":[
"Bergskam",
"bergskrön",
"berg",
"dal",
"dalgång"
],
"natural/sand":[
"Sand",
"strand",
"öken"
],
"natural/scree":[
"röse",
"lösa block",
"stenanhopning",
"Stensamling",
"block",
"stenras",
"Taluskon"
],
"natural/scrub":[
"busksnår",
"sly",
"Buskskog",
"snår"
],
"natural/spring":[
"källsprång",
"springflöde",
"Källa",
"källåder",
"källa",
"vattenställe",
"källdrag",
"källflöde",
"vattenhål"
],
"natural/tree":[
"lövträd",
"ek",
"trä",
"träd",
"barrträd",
"gran",
"Träd",
"stam",
"stock",
"trädstam",
"björk"
],
"natural/tree_row":[
"Träallé",
"trädrad",
"boulevard",
"allé",
"aveny",
"trädkantad väg",
"Trädrad",
"lövgång",
"esplanad"
],
"natural/volcano":[
"lava",
"berg",
"vulkankrater",
"magma",
"krater",
"Vulkan"
],
"natural/water":[
"vattensamling",
"damm",
"reservoar",
"Vatten",
"göl",
"tjärn",
"vatten",
"sjö"
],
"natural/water/lake":[
"insjö",
"vattensamling",
"lagun",
"pöl",
"tjärn",
"göl",
"vatten",
"Sjö",
"innanhav"
],
"natural/water/pond":[
"damm",
"kvarndamm",
"Tjärn",
"liten sjö",
"tjärn",
"göl"
],
"natural/water/reservoir":[
"fördämning",
"Reservoar",
"damm",
"reservoar",
"tank"
],
"natural/wetland":[
"Våtmark",
"mad",
"sump",
"moras",
"sankmark",
"myr",
"mosse",
"träsk",
"torvmark",
"kärr",
"sumpmark"
],
"natural/wood":[
"vildmark",
"skog",
"Urskog",
"bush",
"regnskog",
"träd",
"djungel",
"Skog (utan skogsbruk)"
],
"noexit/yes":[
"vägslut",
"Återvändsgata",
"blindgata återvändsgata",
"Återvändsgränd"
],
"office":[
"tjänsteman",
"byrå",
"tjänstemän",
"Kontor",
"expedition",
"tjänster"
],
"office/accountant":[
"bokhållare",
"bokföring",
"tjänsteman",
"Bokhållare",
"kontorist",
"räkenskap",
"Redovisningsekonom"
],
"office/administrative":[
"Lokal myndighet"
],
"office/adoption_agency":[
"adoptering",
"Adoptionsbyrå",
"barnupptagande",
"Adoption",
"adoptera"
],
"office/advertising_agency":[
"Reklambyrå",
"annons",
"annonsbyrå",
"reklam",
"marknadsföring",
"annonsering"
],
"office/architect":[
"ritningar",
"byggnadskonstnär",
"Arkitektbyrå",
"arkitektkontor",
"byggnadskonst",
"Arkitekt"
],
"office/association":[
"Frivilligorganisation",
"ideell",
"förening",
"volontär",
"organisation",
"frivilligarbetare",
"samhälle",
"icke vinstdrivande",
"Frivillig",
"biståndsarbetare"
],
"office/charity":[
"Välgörenhet",
"biståndsorganisation",
"hjälpverksamhet",
"Välgörenhetsorganisation",
"bistånd"
],
"office/company":[
"expedition",
"kontor",
"Företagskontor",
"kundmottagning",
"företag"
],
"office/coworking":[
"distansarbete",
"mötesrum",
"kontor",
"lånekontor",
"Dagkontor",
"affärslounger",
"tillfällig arbetsplats",
"Coworking",
"Kontorsplats",
"kontorsarbetsplats",
"tillfälligt kontor",
"fjärrarbetsplats",
"konferensrum"
],
"office/educational_institution":[
"rektorsexpedition",
"skolledning",
"rektor",
"skolexpedition",
"Utbildningskontor",
"expedition"
],
"office/employment_agency":[
"förmedling",
"Arbetsförmedling",
"arbetsförmedlingen",
"jobb",
"arbetssökande",
"arbetslös"
],
"office/energy_supplier":[
"ström",
"el",
"gas",
"Elbolag",
"Energibolag",
"energi"
],
"office/estate_agent":[
"fastighet",
"husförmedling",
"mäklare",
"Bostadsförmedling",
"fastighetsmäklare",
"fastighetsuthyrning",
"fastighetsförmedling",
"Mäklare/bostadsförmedling",
"egendom",
"bostadsuthyrning",
"mark",
"kontorsuthyrning"
],
"office/financial":[
"finans",
"bank",
"Bankkontor",
"ekonomisk",
"ekonomi",
"finanskontor"
],
"office/forestry":[
"skog",
"Skogsbolag",
"skogsvaktare"
],
"office/foundation":[
"Stiftelse",
"donation",
"fond"
],
"office/government":[
"myndighetskontor",
"statlig myndighet",
"Myndighet"
],
"office/government/register_office":[
"stadshus",
"inskrivningskontor",
"Folkbokföring",
"registreringskontor",
"Skattemyndigheten",
"mantalslängder",
"registrerade enhet",
"Registreringsbyrå",
"borgerlig vigsel"
],
"office/government/tax":[
"Skattekontor",
"skattemyndigheten",
"myndighet",
"skatt"
],
"office/guide":[
"Turistguide",
"Guidekontor",
"Fjällguide",
"Rundtur",
"Dykguide",
"guide"
],
"office/insurance":[
"försäkringar",
"försäkringsförmedling",
"Försäkringskontor"
],
"office/it":[
"mjukvaruutveckling",
"hårdvara",
"it-specialist",
"IT-kontor",
"it",
"datorer",
"program",
"datorspecialist",
"datakonsult",
"konsultkontor",
"programmering",
"datorkonsult",
"dator",
"systemutveckling",
"mjukvara",
"konsult"
],
"office/lawyer":[
"advokat",
"juridiskt ombud",
"jurist",
"lagman",
"rättsombud",
"ombud",
"Advokatkontor",
"försvarare"
],
"office/lawyer/notary":[
"Notariekontor"
],
"office/moving_company":[
"flytt",
"flyttlass",
"Flyttfirma",
"bärare",
"flyttning",
"transport",
"flyttkarl"
],
"office/newspaper":[
"redaktion",
"utgivare",
"nyhetsredaktion",
"tidning",
"Tidningsredaktion",
"tidningslokal",
"magasin",
"tidskrift"
],
"office/ngo":[
"frivillig",
"ideell förening",
"frivilligorganisation",
"intresseorganisation",
"ideell",
"förening",
"icke-kommersiell",
"organisation",
"hjälporganisation",
"fackförening",
"Icke-statlig organisation"
],
"office/notary":[
"Notarie",
"arv",
"avtal",
"värdehandlningar",
"bevittna",
"egendom",
"fullmakt",
"handlingar",
"Notarius",
"testamente",
"namnteckning",
"dödsbo",
"Notariekontor",
"underskrift",
"signatur",
"Notarius publicus",
"kontrakt",
"påskrift"
],
"office/physician":[
"Läkare"
],
"office/political_party":[
"Politiskt parti",
"politik",
"parti"
],
"office/private_investigator":[
"detektiv",
"deckare",
"Privatdetektiv"
],
"office/quango":[
"Kvasiautonom icke-statlig organisation",
"kvasi",
"organisation",
"Kvasiautonom",
"icke-statlig",
"Quango"
],
"office/research":[
"efterforskning",
"undersökning",
"forskning",
"utveckling",
"vetenskapligt studium",
"vetenskapligt arbete",
"Forskning och utveckling",
"research"
],
"office/surveyor":[
"riskbedömare",
"riskbedömning",
"Undersökning",
"Undersökning/inspektion",
"inspektion",
"stickprovsundersökning",
"statistik",
"enkät",
"lantmätare",
"opinionsundersökning",
"skadebedömare",
"skadebedömning",
"lantmäteri",
"mätning"
],
"office/tax_advisor":[
"ekonomirådgivning",
"Skatterådgivning",
"skattekonsultation",
"skatteplanering",
"moms",
"ekonomi",
"konsultation",
"skatt"
],
"office/telecommunication":[
"mobiltelefon",
"mobiltelefoni",
"surfning",
"internetcafé",
"telefoni",
"telefon",
"Telekom",
"telefoner",
"surfcafé mobil",
"internet"
],
"office/therapist":[
"Radioterapi",
"beteendeterapi",
"Psykoterapi",
"Talterapi",
"psykolog",
"Språkterapi",
"Psykoanalys",
"Samtalsterapi",
"psykologi",
"behandling",
"Kognitiv beteendeterapi",
"Arbetsterapi",
"cellgiftsbehandling",
"sjukgymnast",
"Kemoterapi",
"Farmakoterapi",
"Terapeut",
"Familjeterapi",
"behandlare",
"psykoterapeut",
"Röstterapi",
"Beteendeterapi",
"logoped",
"terapi",
"arbetsterapeut",
"Sexterapi",
"Kognitiv terapi",
"Fysioterapi",
"kbt"
],
"office/travel_agent":[
"Resebyrå "
],
"office/water_utility":[
"Dricksvatten",
"Vattenleverantör",
"vattenbolag"
],
"piste/downhill":[
"skidor",
"alpint",
"slalombacke",
"Utförsåkning",
"skidbacke",
"pist",
"snowboard"
],
"piste/hike":[
"vintervandring",
"vandring",
"snöskor",
"skidor",
"Snöskorvandring",
"vandringsled",
"Snöskorvandring eller vintervandring",
"pist"
],
"piste/ice_skate":[
"isbana",
"skridskor",
"skridskoåkning",
"Skridskoled",
"skridskobana",
"is",
"pist"
],
"piste/nordic":[
"Längdskidåkning eller off-pist/Skidspår",
"off-pist",
"skidor",
"Längdskidåkning",
"skating",
"skidspår",
"pist",
"längdskidor"
],
"piste/piste":[
"isåkning",
"off-pist",
"vintervandring",
"skridsko",
"skidor",
"utför",
"skidtur",
"släde",
"Vintersportspår",
"alpint",
"skida",
"is",
"utförsåkning",
"häst",
"skidåkning",
"snöskor",
"skridskoåkning",
"offpist",
"snowboard"
],
"piste/skitour":[
"skidturåkning",
"skidåkning",
"skidtur",
"skidor",
"skidspår",
"Skidturspår",
"pist"
],
"piste/sled":[
"skidor",
"släde",
"Slädspår",
"slädpist",
"pist"
],
"piste/sleigh":[
"skidor",
"släde",
"Slädspår",
"slädpist",
"pist"
],
"place":[
"Plats"
],
"place/city":[
"stad",
"metropol",
"storstad",
"världsstad",
"huvudstad",
"Större stad"
],
"place/city_block":[
"bostadskomplex",
"husgrupp",
"Kvarter"
],
"place/farm":[
"Gård"
],
"place/hamlet":[
"småort",
"gårdar",
"By",
"litet samhälle",
"gårdssamling"
],
"place/island":[
"holme",
"klippa",
"atoll",
"rev",
"skär",
"ö",
"kobbe",
"Ö",
"skärgård"
],
"place/islet":[
"holme",
"atoll",
"grynna",
"grund",
"rev",
"skär",
"ö",
"kobbe",
"liten ö",
"Holme",
"havsklippa",
"skärgård"
],
"place/isolated_dwelling":[
"bosättning",
"Isolerad boplats",
"boplats"
],
"place/locality":[
"läge",
"lokalitet",
"ställe",
"trakt",
"Plats",
"obefolkad plats"
],
"place/neighbourhood":[
"bostadsområde",
"område",
"närområde",
"stadsdel",
"Kvarter"
],
"place/plot":[
"lott",
"hustomt",
"tomt",
"privat",
"skifte",
"Tomt",
"trädgård",
"mark"
],
"place/quarter":[
"Kvarter / Under-Borough",
"område",
"Under-Borough",
"grannskap",
"stadsdel",
"Kvarter"
],
"place/square":[
"plaza",
"salutorg",
"marknadsplats",
"torg",
"Torg",
"publik yta",
"stadstorg"
],
"place/suburb":[
"kranskommun",
"förort",
"kommundelsnämnd",
"Borough",
"område",
"stadsområde",
"Förort / Borough",
"förstad",
"kommun",
"grannskap",
"stadsdel"
],
"place/town":[
"ort",
"stad",
"Mellanstor stad",
"samhälle"
],
"place/village":[
"ort",
"tätort",
"Mindre samhälle"
],
"playground/balance_beam":[
"Balansbom (lekplats)",
"bom",
"lek",
"lekplats",
"lekområde",
"balansbom",
"balans",
"lekpark"
],
"playground/basket_spinner":[
"karusell",
"lek",
"lekplats",
"lekområde",
"lekpark",
"Korgkarusell"
],
"playground/basket_swing":[
"lek",
"lekplats",
"lekområde",
"gunga",
"kompisgunga",
"Korggunga",
"korg",
"fågelbogunga",
"gungställning",
"lekpark"
],
"playground/climbing_frame":[
"Klätterställning",
"klättring",
"lek",
"lekplats",
"lekområde",
"klättra",
"lekpark"
],
"playground/cushion":[
"Hoppkudde",
"lek",
"lekplats",
"lekområde",
"hoppkudde",
"lekpark"
],
"playground/horizontal_bar":[
"bar",
"lek",
"lekplats",
"lekområde",
"räck",
"lekpark",
"Räck (lekplats)"
],
"playground/rocker":[
"Fjädergunga",
"lek",
"lekplats",
"lekområde",
"Gungdjur",
"lekpark"
],
"playground/roundabout":[
"karusell",
"lek",
"lekplats",
"lekområde",
"Karusell (lekplats)",
"lekpark"
],
"playground/sandpit":[
"sand",
"Sandlåda",
"lek",
"sandlåda",
"lekplats",
"lekområde",
"lekpark"
],
"playground/seesaw":[
"lek",
"gungbräda",
"lekplats",
"lekområde",
"Gungbräda",
"lekpark"
],
"playground/slide":[
"lek",
"lekplats",
"lekområde",
"Rutschkana",
"rutschbana",
"lekpark",
"rutchelbana"
],
"playground/structure":[
"lek",
"lekplats",
"lekområde",
"Lekhus",
"Lekslott",
"lekhus",
"lekstuga",
"lekpark"
],
"playground/swing":[
"lek",
"Gunga",
"lekplats",
"lekområde",
"Gungställning",
"lekpark"
],
"playground/zipwire":[
"lek",
"lekplats",
"lekområde",
"Linbana (lekplats)",
"linbana",
"lekpark"
],
"point":[
"läge",
"fläck",
"plats",
"ställe",
"Punkt"
],
"power":[
"Elförsörjning"
],
"power/cable/underground":[
"kraft",
"ström",
"högspänning",
"underjordisk kraftkabel",
"Kraftledning",
"elledning",
"elnät",
"El",
"högspänningsledning",
"strömförsörjning",
"elförsörjning",
"Underjordisk kraftkabel"
],
"power/generator":[
"strömtillverkning",
"Elgenerator",
"kraftgenerator",
"kraftkälla",
"generator"
],
"power/generator/method/photovoltaic":[
"solenergi",
"PV-modul",
"fotovoltaik",
"solcell",
"solkraft",
"solljus",
"solkraftverk",
"Solpanel",
"termisk solkraft",
"solcellsmodul",
"solel"
],
"power/generator/source/nuclear":[
"kärnanläggning",
"kärnenergi",
"kärnreaktor",
"atomkraftverk",
"kärnkraft",
"kärnkraftvärk",
"reaktor",
"atomkraft",
"Kärnkraftsreaktor",
"nukleär energi",
"kärnkraftverk",
"atomenergi",
"kärnkraftsanläggning"
],
"power/generator/source/wind":[
"vindmölla",
"Vindturbin",
"vindkraftverk",
"vindkraft"
],
"power/line":[
"kraftledning",
"högspänning",
"elledning",
"högspänningsledning",
"Högspänningsledning"
],
"power/minor_line":[
"Kraftledning",
"elledning",
"Mindre kraftledning"
],
"power/plant":[
"el",
"Kol",
"generator",
"kraft",
"vind*",
"elkraftverk",
"vattenkraft*",
"kärnkraft*",
"Område för kraftproduktion",
"elproduktion",
"gas",
"solkraft*",
"kraftproduktion"
],
"power/pole":[
"elledningsstolpe",
"mast",
"stolpe",
"Kraftledningsstolpe",
"kraftledningsmast",
"elledningsmast"
],
"power/sub_station":[
"Fördelningsstation"
],
"power/substation":[
"elomvandling",
"Fördelningsstation",
"fördelningsstation",
"stadsnätstation",
"elskåp",
"Transformator",
"elfördelning"
],
"power/switch":[
"Strömbrytare",
"Frånskiljare"
],
"power/tower":[
"mast",
"Högspänningsmast",
"kraftledningsstolpe",
"kraftledningsmast"
],
"power/transformer":[
"elomvandling",
"nätstation",
"Transformator"
],
"public_transport/linear_platform":[
"Hållplats",
"kollektivtrafik",
"Plattform",
"linjetrafik",
"transport",
"Hållplats / Plattform för kollektivtrafik"
],
"public_transport/linear_platform_aerialway":[
"linbanestopp",
"hållplats",
"stopp",
"Hållplats / Plattform för linbana",
"linbaneterminal",
"aerialway",
"linbana",
"terminal",
"linjetrafik",
"transport",
"Linbanehållplats",
"kollektivtrafik",
"transit",
"plattform",
"linbaneplattform"
],
"public_transport/linear_platform_bus":[
"busshållplats",
"kollektivtrafik",
"hållplats",
"bussplattform",
"Bussplattform",
"transit",
"plattform",
"transport",
"linjetrafik",
"buss"
],
"public_transport/linear_platform_ferry":[
"brygga",
"stopp",
"båthållplats",
"Färjeterminal",
"Färjestation",
"färjestopp",
"terminal",
"linjetrafik",
"transport",
"färja",
"båt",
"färjeplattform",
"kollektivtrafik",
"båtterminal",
"transit",
"pir",
"station",
"plattform",
"Färjehållplats",
"Stop / plattform för färja",
"båtstopp"
],
"public_transport/linear_platform_light_rail":[
"Hållplats för snabbspårväg / stadsbana",
"hållplats",
"light rail",
"spårvagnsplattform",
"vagn",
"stadsbana",
"terminal",
"transport",
"Spårvägshållplats",
"snabbspårväg",
"spårväg",
"kollektivtrafik",
"spårvagnsterminal",
"transit",
"spårvagn",
"plattform",
"järnväg",
"spår"
],
"public_transport/linear_platform_monorail":[
"monorailstopp",
"stopp",
"Stopp / plattform för monorail",
"enskensbana",
"linjetrafik",
"transport",
"räls",
"monorail",
"monorailplattform",
"kollektivtrafik",
"plattform",
"balkbana",
"spår"
],
"public_transport/linear_platform_subway":[
"Tunnelbaneplattform",
"Tunnelbanestopp / -plattform",
"kollektivtrafik",
"metro",
"plattform",
"Tunnelbanestopp",
"transport",
"tunnelbana",
"järnväg",
"spår",
"underjordisk"
],
"public_transport/linear_platform_train":[
"järnvägsperrong",
"stopp",
"järnvägsplattform",
"linjetrafik",
"transport",
"Järnvägsstopp / -perrong",
"Perrong",
"kollektivtrafik",
"transit",
"tåg",
"plattform",
"Tågstopp",
"järnväg",
"spår"
],
"public_transport/linear_platform_tram":[
"hållplats",
"spårvagnsplattform",
"vagn",
"Spårvagnshållplats / -plattform",
"terminal",
"transport",
"Spårvägshållplats",
"spårväg",
"kollektivtrafik",
"spårvagnsterminal",
"transit",
"spårvagn",
"plattform",
"spårvagnshållplats",
"järnväg"
],
"public_transport/linear_platform_trolleybus":[
"Busshållplats",
"hållplats",
"spårlös",
"vagn",
"transport",
"trådbuss",
"kollektivtrafik",
"bussplattform",
"transit",
"spårvagn",
"Busshållplats / plattform för trådbuss",
"plattform",
"buss"
],
"public_transport/platform":[
"väntplats",
"avsats",
"Plattform",
"påstigningsplats",
"perrong",
"Stopp / Plattform för kollektivtrafik"
],
"public_transport/platform_aerialway":[
"linbanestopp",
"hållplats",
"stopp",
"Hållplats / Plattform för linbana",
"linbaneterminal",
"aerialway",
"linbana",
"terminal",
"linjetrafik",
"transport",
"Linbanehållplats",
"kollektivtrafik",
"transit",
"plattform",
"linbaneplattform"
],
"public_transport/platform_bus":[
"busshållplats",
"kollektivtrafik",
"hållplats",
"bussplattform",
"transit",
"plattform",
"transport",
"linjetrafik",
"Busshållplats / Bussplattform",
"buss"
],
"public_transport/platform_ferry":[
"brygga",
"stopp",
"båthållplats",
"Färjeterminal",
"Färjestation",
"färjestopp",
"terminal",
"linjetrafik",
"transport",
"färja",
"båt",
"färjeplattform",
"kollektivtrafik",
"båtterminal",
"transit",
"pir",
"station",
"plattform",
"Färjehållplats",
"Stop / plattform för färja",
"båtstopp"
],
"public_transport/platform_light_rail":[
"Hållplats för snabbspårväg / stadsbana",
"hållplats",
"light rail",
"spårvagnsplattform",
"vagn",
"stadsbana",
"terminal",
"transport",
"Spårvägshållplats",
"snabbspårväg",
"spårväg",
"kollektivtrafik",
"spårvagnsterminal",
"transit",
"spårvagn",
"plattform",
"järnväg",
"spår"
],
"public_transport/platform_monorail":[
"monorailstopp",
"stopp",
"Stopp / plattform för monorail",
"enskensbana",
"linjetrafik",
"transport",
"räls",
"monorail",
"monorailplattform",
"kollektivtrafik",
"plattform",
"balkbana",
"spår"
],
"public_transport/platform_subway":[
"Tunnelbaneplattform",
"Tunnelbanestopp / -plattform",
"kollektivtrafik",
"metro",
"plattform",
"Tunnelbanestopp",
"transport",
"tunnelbana",
"järnväg",
"spår",
"underjordisk"
],
"public_transport/platform_train":[
"järnvägsperrong",
"stopp",
"järnvägsplattform",
"linjetrafik",
"transport",
"Järnvägsstopp / -perrong",
"Perrong",
"kollektivtrafik",
"transit",
"tåg",
"plattform",
"Tågstopp",
"järnväg",
"spår"
],
"public_transport/platform_tram":[
"hållplats",
"spårvagnsplattform",
"vagn",
"Spårvagnshållplats / -plattform",
"terminal",
"transport",
"Spårvägshållplats",
"spårväg",
"kollektivtrafik",
"spårvagnsterminal",
"transit",
"spårvagn",
"plattform",
"spårvagnshållplats",
"järnväg"
],
"public_transport/platform_trolleybus":[
"Busshållplats",
"hållplats",
"spårlös",
"vagn",
"transport",
"trådbuss",
"kollektivtrafik",
"bussplattform",
"transit",
"spårvagn",
"Busshållplats / plattform för trådbuss",
"plattform",
"buss"
],
"public_transport/station":[
"kollektivtrafik",
"Station för kollektivtrafik",
"bytespunkt",
"station",
"resecenter",
"terminal",
"transport"
],
"public_transport/station_aerialway":[
"kollektivtrafik",
"transit",
"Linbanestation",
"station",
"aerialway",
"linbana",
"terminal",
"transport"
],
"public_transport/station_bus":[
"Busshållplats",
"kollektivtrafik",
"transit",
"station",
"resecenter",
"Bussterminal",
"reseterminal",
"terminal",
"transport",
"Busstation / Bussterminal",
"Busstation",
"buss"
],
"public_transport/station_ferry":[
"brygga",
"Färjeterminal",
"båthållplats",
"Färjestation",
"terminal",
"transport",
"färja",
"båt",
"kollektivtrafik",
"Färjeterminal / Färjehållplats / Färjestation",
"båtterminal",
"transit",
"pir",
"station",
"Färjehållplats"
],
"public_transport/station_light_rail":[
"light rail",
"lättbana",
"hållplats",
"stadsbana",
"spårvagnstopp",
"Station för snabbspårväg / stadsbana",
"transport",
"linjetrafik",
"terminal",
"snabbspårväg",
"spårväg",
"kollektivtrafik",
"spårvagnsterminal",
"Station för snabbspårväg",
"spårvagn",
"station",
"spårvagnshållplats",
"Station för light rail",
"järnväg",
"spår"
],
"public_transport/station_monorail":[
"enskensbana",
"terminal",
"linjetrafik",
"transport",
"monorailstation",
"räls",
"monorail",
"kollektivtrafik",
"station",
"plattform",
"Monorailstation",
"spår",
"balkbana"
],
"public_transport/station_subway":[
"",
"kollektivtrafik",
"metro",
"station",
"transport",
"terminal",
"tunnelbana",
"järnväg",
"spår",
"underjordisk",
"Tunnelbanestation"
],
"public_transport/station_train":[
"linjeplats",
"trafikplats",
"central",
"tåghållplats",
"hållplats",
"Järnvägsstation",
"järnvägshållplats",
"centralstation",
"huvudbangård",
"hållställe",
"tågstation"
],
"public_transport/station_train_halt":[
"hållplats",
"hållställe",
"transport",
"avstigning",
"Mindre järnvägshållplats",
"kollektivtrafik",
"järnvägshållplats",
"påstigning",
"transit",
"tåg",
"station",
"plattform",
"järnvägsstation",
"järnväg",
"spår"
],
"public_transport/station_tram":[
"spårväg",
"Spårvagnsstation",
"spårvagnsterminal",
"spårvagn",
"station",
"spårvägshållplats"
],
"public_transport/station_trolleybus":[
"busshållplats",
"hållplats",
"terminal",
"linjetrafik",
"transport",
"Station / Terminal för trådbuss",
"trådbussterminal",
"trådbuss",
"trådbusstopp",
"kollektivtrafik",
"bussterminal",
"station",
"busstopp",
"trådbusshållplats",
"buss"
],
"public_transport/stop_area":[
"kollektivtrafik",
"hållplats",
"bytespunkt",
"transit",
"byte",
"station",
"knutpunkt",
"resecenter",
"terminal",
"linjetrafik",
"transport",
"Bytespunkt / knutpunkt"
],
"public_transport/stop_position":[
"stopposition",
"kollektivtrafik",
"hållplats",
"Stopposition för kollektivtrafik",
"linjetrafik",
"transport"
],
"public_transport/stop_position_aerialway":[
"Stopposition för linbana",
"stopposition",
"linbanestation",
"linbanestopp",
"kollektivtrafik",
"hållplats",
"linbaneterminal",
"linbana",
"linjetrafik",
"transport",
"linbanehållplats"
],
"public_transport/stop_position_bus":[
"stopposition",
"busshållplats",
"kollektivtrafik",
"hållplats",
"bussterminal",
"busstopp",
"linjetrafik",
"transport",
"buss",
"Stopposition för buss"
],
"public_transport/stop_position_ferry":[
"båt",
"stopposition",
"busshållplats",
"kollektivtrafik",
"hållplats",
"bussterminal",
"busstopp",
"linjetrafik",
"transport",
"Stopposition för färja",
"färja"
],
"public_transport/stop_position_light_rail":[
"stopposition",
"light rail",
"lättbana",
"hållplats",
"stadsbana",
"spårvagnstopp",
"transport",
"linjetrafik",
"snabbspårväg",
"spårväg",
"kollektivtrafik",
"spårvagnsterminal",
"spårvagn",
"Stopposition för snabbspårväg / stadsbana",
"spårvagnshållplats",
"Stopposition för snabbspårväg",
"järnväg",
"spår"
],
"public_transport/stop_position_monorail":[
"stopposition",
"kollektivtrafik",
"hållplats",
"Stopposition för monorail",
"enskensbana",
"linjetrafik",
"transport",
"balkbana",
"spår",
"räls",
"monorail"
],
"public_transport/stop_position_subway":[
"tunnelbanetåg",
"stopposition",
"tunnelbanestation",
"kollektivtrafik",
"hållplats",
"tunnelbanestopp",
"linjetrafik",
"transport",
"tunnelbana",
"tunnelbanehållplats",
"Stopposition för tunnelbana"
],
"public_transport/stop_position_train":[
"tågterminal",
"järnvägsstopp",
"stopposition",
"hållplats",
"linjetrafik",
"transport",
"tågstopp",
"kollektivtrafik",
"järnvägshållplats",
"tåg",
"järnvägsterminal",
"järnvägsstation",
"Stopposition för tåg",
"tågstation"
],
"public_transport/stop_position_tram":[
"stopposition",
"kollektivtrafik",
"hållplats",
"spårvagnsterminal",
"Stopposition för spårvagn",
"spårvagn",
"spårvagnstopp",
"spårvagnshållplats",
"linjetrafik",
"transport"
],
"public_transport/stop_position_trolleybus":[
"stopposition",
"busshållplats",
"hållplats",
"Stopposition för trådbuss",
"linjetrafik",
"transport",
"trådbussterminal",
"trådbuss",
"trådbusstopp",
"kollektivtrafik",
"bussterminal",
"busstopp",
"trådbusshållplats",
"buss"
],
"railway":[
"Järnväg"
],
"railway/abandoned":[
"borttagen järnväg",
"Riven järnväg"
],
"railway/buffer_stop":[
"Stoppbock",
"Buffertstopp",
"Buffert",
"stoppblock"
],
"railway/crossing":[
"spårpassage",
"järnvägspassage",
"cykelväg",
"gångväg",
"stig",
"tågkorsning",
"plankorsning",
"tågövergång",
"cykelpassage",
"Järnvägskorsning (stig)",
"gångpassage",
"järnvägskorsning",
"tågpassage",
"korsning",
"järnvägsövergång",
"övergångsställe"
],
"railway/derail":[
"utspårare",
"Spårspärr",
"omläggningsanordning"
],
"railway/disused":[
"övergiven järnväg",
"oanvänd tågbana",
"övergiven tågbana",
"Oanvänd järnväg"
],
"railway/funicular":[
"Bergbana ",
"linbana",
"Bergbana"
],
"railway/halt":[
"Mindre järnvägshållplats"
],
"railway/level_crossing":[
"spårpassage",
"järnvägspassage",
"tågkorsning",
"plankorsning",
"tågövergång",
"järnvägskorsning",
"Järnvägskorsning (väg)",
"tågpassage",
"korsning",
"järnvägsövergång"
],
"railway/light_rail":[
"smalspår",
"smalspårig järnväg",
"Snabbspårväg / stadsbana",
"stadsbana",
"järnväg",
"snabbspårväg"
],
"railway/milestone":[
"Kilometerstolpe",
"kilometertavla",
"kilometerpåle",
"milsten",
"referenstavla",
"Kilometerstolpe vid järnväg",
"avståndsmärke"
],
"railway/miniature":[
"smalspår",
"smalspårig järnväg",
"trädgårdsjärnväg",
"Åkbar miniatyrjärnväg",
"Miniatyrjärnväg"
],
"railway/monorail":[
"Monorail",
"kollektivtrafik",
"enskensbana",
"linjetrafik",
"transport",
"balkbana",
"spår",
"räls"
],
"railway/narrow_gauge":[
"smalspår",
"Smalspårbana"
],
"railway/platform":[
"Järnvägsstopp / -perrong"
],
"railway/rail":[
"Räls",
"järnvägsspår",
"spår",
"bana"
],
"railway/signal":[
"semafor",
"huvudsignal",
"järnvägssignal",
"järnvägsljus",
"försignal",
"signal",
"ljus",
"Järnvägssignal",
"dvärgsignal"
],
"railway/station":[
"Järnvägsstation"
],
"railway/subway":[
"T-bana",
"metro",
"Tunnelbana"
],
"railway/subway_entrance":[
"Tunnelbaneingång",
"t-banenedgång",
"t-baneingång",
"tunnelbanenergång"
],
"railway/switch":[
"korsningsväxel",
"järnvägskorsning",
"växel",
"Järnvägsväxel",
"korsning"
],
"railway/train_wash":[
"tvätthall",
"Tågtvätt",
"loktvätt"
],
"railway/tram":[
"Spårvagn",
"spårväg",
"motorvagn"
],
"railway/tram_stop":[
"Stopposition för spårvagn"
],
"relation":[
"Relation",
"samband",
"relaterat",
"koppling",
"anknytning",
"förbindelse",
"förhållande",
"kontext"
],
"roundabout":[
"Cirkulationsplats"
],
"route/ferry":[
"färjelinje",
"båtlinje",
"båtrutt",
"rutt",
"Färjerutt",
"färja",
"båt i linjetrafik"
],
"seamark":[
"Sjöfart"
],
"shop":[
"shop",
"butik",
"Affär"
],
"shop/agrarian":[
"utsäde",
"jordbruksmaskiner",
"frön",
"Jordbruksaffär",
"gödsel",
"djurmat",
"gödningsmedel",
"jordbruksverktyg",
"lantmannaföreningen",
"bekämpningsmedel",
"jordbruksutrustning",
"Jordbruk"
],
"shop/alcohol":[
"spritaffär",
"systemet",
"öl",
"systembolaget",
"Vin-och-spritaffär",
"bolaget",
"vin- och spritaffär",
"alkohol",
"sprit",
"vin- och sprit",
"vin",
"Vinaffär"
],
"shop/anime":[
"animēshon",
"Anime-affär",
"Anime",
"Josei",
"Kodomo",
"Shōjo",
"manga",
"mangastil",
"shojo",
"shoujo",
"Shōnen"
],
"shop/antiques":[
"antikvitetsaffär",
"antikt",
"Antikaffär",
"antikshop",
"antikvariat"
],
"shop/appliance":[
"tvättmaskin",
"vitvarukedja",
"vitvaruaffär",
"mikrovågsugn",
"köksfläkt",
"spis",
"frys",
"hushållsmaskin",
"Vitvaror",
"hushållsmaskiner",
"kylskåp",
"ugn",
"vitvaror",
"vitvara",
"diskmaskin"
],
"shop/art":[
"konstverk",
"Konstaffär",
"tavlor",
"kulturer",
"konst",
"konsthandlare",
"konstgalleri",
"galleri",
"statyer",
"konstutställning"
],
"shop/baby_goods":[
"Bäbis",
"Babyprodukter",
"småbarn",
"nappflaskor",
"nappar",
"babykläder",
"Baby",
"barnkläder",
"bäbiskläder",
"barnvagnar",
"spjälsängar",
"blöjor"
],
"shop/bag":[
"bagageväskor",
"resväskor",
"bagage",
"handväska",
"väskor",
"Väskaffär",
"plånbok",
"handväskor"
],
"shop/bakery":[
"bröd",
"Bageri",
"bullar",
"baka",
"bagare"
],
"shop/bathroom_furnishing":[
"Badrumsinredning",
"badrum"
],
"shop/beauty":[
"Skönhetssalong",
"nagelsalong",
"spa",
"skönhet",
"kuranstalt",
"smink",
"salong",
"kosmetik",
"solarium",
"shiatsu",
"hälsoanläggning",
"kurort",
"naglar",
"skönhetsbehandlingar",
"massage"
],
"shop/beauty/nails":[
"nagel",
"nagelvård",
"naglar",
"manikur",
"handvård",
"händer",
"manikyr",
"Nagelsalong",
"pedikyr",
"hand",
"manikyrist  manikyrera"
],
"shop/beauty/tanning":[
"solarium",
"konstgjort solljus",
"Solarium"
],
"shop/bed":[
"madrasser",
"Sängaffär",
"sängar",
"påslakan",
"täcken",
"lakan",
"kuddar"
],
"shop/beverages":[
"Dryck",
"dricka",
"läsk",
"alkohol",
"Dryckaffär",
"läskedryck"
],
"shop/bicycle":[
"cykelförsäljning",
"Cykelaffär",
"cykel",
"cykelreparatör"
],
"shop/bookmaker":[
"spel",
"Stryktipset",
"måltipset",
"trav",
"Vadslagning",
"dobbel",
"vadhållning"
],
"shop/books":[
"Bokhandel",
"antikvariat",
"bokförsäljning"
],
"shop/boutique":[
"smycken",
"Boutique (Dyra kläder och accessoarer)",
"finkläder",
"Boutique",
"modeaffär",
"accessoarer",
"klänningar",
"kläder"
],
"shop/butcher":[
"Slaktare",
"köttaffär",
"charkuterihandlare",
"chark",
"köttstyckare",
"slaktare",
"styckare",
"kött",
"charkuterist"
],
"shop/candles":[
"värmeljus",
"Ljusaffär",
"mysljus",
"ljusstakar",
"ljus",
"stearinljus"
],
"shop/car":[
"bilfirma",
"bilreparatör",
"bilförsäljning",
"bilverkstad",
"bilsäljare",
"Bilhandlare",
"biltillbehör"
],
"shop/car_parts":[
"Bildelar",
"bilreservdelar",
"motor",
"Biltillbehör",
"reservdelar",
"biltillbehör"
],
"shop/car_repair":[
"motor",
"bilreparatör",
"Bilverkstad",
"verkstad"
],
"shop/carpet":[
"matta",
"Mattaffär",
"mattor"
],
"shop/charity":[
"myrorna",
"begagnat",
"secondhandbutik",
"välgörenhetsbutik",
"andrahandsbutik",
"second hand",
"secondhand",
"second hand-butik",
"begagnade varor",
"bättre begagnat",
"vintage",
"Second hand-butik",
"second handbutik",
"välgörenhet"
],
"shop/cheese":[
"ost",
"ostar",
"Ostaffär",
"ostbutik"
],
"shop/chemist":[
"hygienartiklar",
"kosmetik",
"kemi",
"Kemiaffär",
"städ",
"rengöring",
"smink",
"hygien",
"kosmetika",
"städmaterial",
"Kemiaffär (hygien,  kosmetika & städ)",
"rengöringsmedel"
],
"shop/chocolate":[
"pralin",
"konfekt",
"Chokladaffär",
"Choklad",
"praliner"
],
"shop/clothes":[
"klädbutik",
"ekipering",
"Klädaffär",
"kläder"
],
"shop/coffee":[
"kaffeaffär",
"kaffepulver",
"Kaffeaffär",
"kaffeböner",
"kaffebönor",
"bryggkaffe",
"kaffe"
],
"shop/computer":[
"data",
"dator",
"datorförsäljning",
"Datorbutik",
"datorer",
"datoraffär",
"datorhårdvara",
"datorprogram"
],
"shop/confectionery":[
"konfektyr",
"choklad",
"sötsaker",
"godisbutik",
"godisaffär",
"godis",
"Godisaffär",
"konfektbutik",
"karameller"
],
"shop/convenience":[
"livsmedelsbutik",
"mataffär",
"Närbutik",
"kvartersbutik",
"livsmedel"
],
"shop/copyshop":[
"kopiering",
"Tryckeri",
"tryckeri",
"Copyshop"
],
"shop/cosmetics":[
"Sminkaffär",
"smink",
"kosmetika",
"kosmetikaffär"
],
"shop/craft":[
"konstverk",
"hantverk",
"Konsthantverk",
"slöjd",
"Konst- och hantverksbutik"
],
"shop/curtain":[
"Gardinaffär",
"drapera",
"fönster",
"draperier",
"gardiner"
],
"shop/dairy":[
"ost",
"ägg",
"mejeri",
"mjölk",
"mjölkaffär",
"Mejeriaffär"
],
"shop/deli":[
"lunch",
"smörgås",
"delikatess",
"Delikatessaffär",
"delikatesser",
"finmat",
"kött"
],
"shop/department_store":[
"Varuhus",
"affärshus"
],
"shop/doityourself":[
"indie",
"handverktyg",
"heminredning",
"elverktyg",
"byggvaruhus",
"inredning",
"byggsatser",
"verktyg",
"byggsats",
"Gör-det-själv",
"gördetsjälv",
"gör det själv",
"Byggmarknad",
"byggmaterial",
"järnaffär",
"bygghandel"
],
"shop/dry_cleaning":[
"Kemtvättar",
"Kemtvätt",
"kemisk tvätt"
],
"shop/e-cigarette":[
"elektrisk cigarett",
"elcigarett",
"Affär för elektroniska cigaretter",
"e-cigarett"
],
"shop/electronics":[
"spisar",
"TV",
"batterier",
"tvättmaskin",
"kablar",
"datorer",
"radio",
"apparater",
"dator",
"hemelektronik",
"kylskåp",
"torktumlare",
"Elektronikbutik",
"vitvaror",
"hushållsapparater",
"ljud"
],
"shop/erotic":[
"erotik",
"sexaffär",
"Sex",
"sexleksaker",
"sexshop",
"porr",
"pornografi",
"porrfilmer",
"Sexshop",
"erotikaffär",
"porrtidningar",
"underkläder",
"sexfilmer",
"kondomer",
"erotisk"
],
"shop/fabric":[
"Tygaffär",
"tyg",
"tyger",
"sy",
"sömnad"
],
"shop/farm":[
"närproducerat",
"Gårdsbutik",
"egenproducerat"
],
"shop/fashion":[
"mode",
"Modebutik",
"modekläder",
"klädaffär",
"kläder"
],
"shop/fishmonger":[
"Fiskhandlare"
],
"shop/florist":[
"Florist",
"bukett",
"blomsterhandlare",
"blommor",
"blomsterbindare",
"blomförsäljning"
],
"shop/frame":[
"Ramaffär",
"ramar",
"inramning"
],
"shop/funeral_directors":[
"gravsten",
"bodelning",
"begravning",
"jordfästning",
"gravsättning",
"begravningsentreprenör",
"Begravningsbyrå",
"kremering",
"begravningsbyrå",
"gravstenar",
"begravningsceremoni"
],
"shop/furnace":[
"Värmepannor"
],
"shop/furniture":[
"möbelgrossist",
"bord",
"hylla",
"soffor",
"inredning",
"stol",
"Möbelaffär",
"stolar",
"möbelvaruhus",
"soffa"
],
"shop/garden_centre":[
"krukväxter",
"trädgårdsväxter",
"jord",
"Trädgårdscenter",
"träd",
"trädgårdsverktyg",
"planteringsjord",
"kompost",
"blomkrukor",
"blommor",
"landskap",
"plantskola",
"buskar",
"trädgård"
],
"shop/gas":[
"gasbehållare",
"lpg",
"metangas",
"gasflaskor",
"propan",
"Försäljning av gas",
"naturgas",
"gasol",
"fordonsgas",
"återfyllning",
"gas",
"cng",
"gasolflaskor"
],
"shop/gift":[
"gratulationskort",
"souvenirbutik",
"grattiskort",
"presenter",
"souvenirer",
"gåva",
"present",
"Presentbutik",
"gåvor",
"souvenir"
],
"shop/greengrocer":[
"frukt",
"frukthandlare",
"grönsaker",
"frukthandel",
"Grönsakshandlare",
"vegetabiliskt"
],
"shop/hairdresser":[
"hårkonstnär",
"skägg",
"skönhet",
"skönhetssalong",
"hårförlängning",
"hårkreatör",
"salong",
"stylist",
"hårklippning",
"barberare",
"rakning",
"frisör",
"hår",
"hårtvätt",
"hårfärgning",
"Hårfrisör"
],
"shop/hardware":[
"handverktyg",
"nycklar",
"spik",
"järntillbehör",
"hushållsprodukter",
"redskap",
"Järnaffär",
"metallverktyg",
"bultar",
"bygg",
"lås",
"kök",
"elverktyg",
"badrum",
"krokar",
"el",
"verktyg",
"skruvar",
"trädgårdsredskap",
"nyckeltillverkning",
"vvs",
"järnhandlare",
"bult",
"järnbeslag",
"köksutrustning",
"skruv"
],
"shop/health_food":[
"Hälsokostbutik",
"kosttillskott",
"hälsokost",
"naturligt",
"organisk",
"köttersättning",
"vegetarian",
"vegan",
"mjölkersättning",
"hälsomat",
"organist",
"vitaminer"
],
"shop/hearing_aids":[
"hörselskada",
"Hörapparater",
"hörselskadade",
"hörsel",
"hörhjälpmedel"
],
"shop/herbalist":[
"läkande örter",
"örter",
"medicinalväxter",
"Medicinalväxter"
],
"shop/hifi":[
"HIFI-butik",
"ljudåtergivning",
"hifi",
"förstärkare",
"stereoanläggning",
"högtalare",
"HiFi-butik",
"ljudanläggning",
"stereo",
"audio",
"video",
"ljud"
],
"shop/houseware":[
"porslin",
"hem",
"köksredskap",
"hushåll",
"husgeråd",
"bestick",
"prydnadsföremål",
"Husgeråd"
],
"shop/interior_decoration":[
"Inredningsaffär",
"inredning",
"dekoration"
],
"shop/jewelry":[
"pärla",
"ringar",
"Juvelerare",
"ring",
"klockor",
"pärlor",
"halsband",
"diamant",
"smycken",
"guld",
"klocka",
"örhängen",
"silver",
"örhänge"
],
"shop/kiosk":[
"glass",
"gatukök",
"läsk",
"dryck",
"tobak",
"tidningar",
"snus",
"snabbmat",
"butik",
"godis",
"korv",
"Kiosk",
"cigaretter"
],
"shop/kitchen":[
"kök",
"bänkskivor",
"köksskåp",
"skåpluckor",
"Köksinredning"
],
"shop/laundry":[
"Tvättinrättning",
"tvättstuga",
"tvättemat",
"tvättautomat",
"tvätteri"
],
"shop/leather":[
"läder",
"läderjackor",
"läderkläder",
"Läderaffär"
],
"shop/locksmith":[
"Låsdyrkning",
"dyrkning",
"nyckel",
"nyckelkopiering",
"Låssmed",
"lås",
"låsinstallation",
"nyckeltillverkning"
],
"shop/lottery":[
"lottförsäljningen",
"bingospel",
"Lotteri",
"lottstånd",
"hasardspel",
"hasard",
"lottdragning",
"tombola"
],
"shop/mall":[
"Köpcenter",
"shoppingcentrum",
"köpcentrum",
"köpcenter",
"Varuhus",
"shoppingcenter",
"affärshus"
],
"shop/massage":[
"massagebehandling",
"thaimassage",
"Massage"
],
"shop/medical_supply":[
"medicinsk utrustning",
"rullstol",
"Bandage",
"blodtrycksmätare",
"Glucometer",
"Träningsbollar",
"Ortopedteknik",
"hjälpmedel",
"ledstöd",
"glukometer",
"Kryckor",
"Medicinsk utrustning "
],
"shop/mobile_phone":[
"mobiltelefon",
"Mobiltelefoner",
"mobiltelefoni",
"telefon",
"telefonbutik",
"mobiltelefonbutik"
],
"shop/money_lender":[
"utlåningsinstitution",
"telefonlån",
"mikrolån",
"pantbank",
"Långivare",
"utlåning"
],
"shop/motorcycle":[
"motorcykelbutik",
"motorcyklar",
"Återförsäljare av motorcyklar",
"Motorcykel",
"motorcykeltillbehör",
"motorcykelåterförsäljare"
],
"shop/motorcycle_repair":[
"motorcykelreparatör",
"motorcyklar",
"motorcykel",
"service",
"cykel",
"Motorcykelverkstad",
"moped",
"reparatör",
"motorcykelservice",
"verkstad",
"reparation",
"mopedverkstad"
],
"shop/music":[
"CD",
"Musikaffär",
"CD-affär",
"kassett",
"LP",
"musikbutik",
"skivaffär",
"vinyl",
"skivbutik"
],
"shop/musical_instrument":[
"noter",
"instrument",
"Musikinstrument"
],
"shop/newsagent":[
"pressbyrå",
"tidskrifter",
"Tidningsaffär",
"pressbyrån",
"tidningar",
"kiosk",
"magasin",
"tidningsställ",
"tidningskiosk"
],
"shop/nutrition_supplements":[
"viktminskning",
"hälsoörter",
"Hälsokost",
"hälsoprodukter",
"hälsa",
"mineraler",
"vitaminer"
],
"shop/optician":[
"glasögon",
"ögon",
"synundersökning",
"linser",
"Optiker"
],
"shop/organic":[
"ekologiskt",
"Ekologiska livsmedel",
"miljövänligt"
],
"shop/outdoor":[
"tält",
"camping",
"klätterutrustning",
"vandring",
"klättring",
"vandringsutrustning",
"uteliv",
"Friluftsaffär",
"campingutrustning",
"friluftsliv"
],
"shop/paint":[
"färg",
"Färgbutik",
"målarfärg",
"målning"
],
"shop/pastry":[
"kondis",
"kaffeservering",
"servering",
"fik",
"sockerbagare",
"kafé",
"konditori",
"café",
"finbageri",
"sockerbageri",
"cafe",
"bageri",
"Konditori"
],
"shop/pawnbroker":[
"pant",
"Pantbank",
"pantbelåning",
"pantbanken",
"pantbank",
"pantlånekontor",
"varubelåning"
],
"shop/perfumery":[
"parfymeri",
"Parfymbutik",
"parfym",
"parfymbutik",
"smink",
"kosmetika"
],
"shop/pet":[
"katter",
"katt",
"Djurbutik",
"hundar",
"djurmat",
"djur",
"akvarium",
"hund",
"fisk",
"djurburar",
"husdjur",
"djurtillbehör",
"Djuraffär"
],
"shop/pet_grooming":[
"hund",
"pälsvård",
"hundvård",
"husdjur",
"Pälsvård för husdjur",
"Trimning"
],
"shop/photo":[
"fotoaffär",
"framkallning",
"kameratillbehör",
"Fotoaffär ",
"fotokamera",
"video",
"film",
"konvertering",
"bild",
"fotografi",
"foto",
"kameror",
"filmkamera",
"fotoredigering",
"kamera",
"ram"
],
"shop/pyrotechnics":[
"Fyrverkerier",
"tomtebloss",
"raketer",
"smällare",
"fyrverkerier",
"pyroteknik",
"nyårsraketer"
],
"shop/radiotechnics":[
"elektronikbutik",
"radiotillbehör",
"radiobutik",
"Radio",
"elektronik",
"elektronikkomponenter",
"Radio/Elektronikbutik"
],
"shop/religion":[
"biblar",
"Religiös",
"kyrkobutik",
"psalmböcker",
"Religiös butik",
"religion"
],
"shop/scuba_diving":[
"Dykning",
"Dykarbutik",
"dykutrustning"
],
"shop/seafood":[
"hummer",
"räkor",
"fisk",
"ostron",
"bläckfisk",
"krabba",
"skaldjur",
"fiskhandlare",
"Fiskaffär",
"musslor"
],
"shop/second_hand":[
"loppis",
"Second hand",
"loppmarknad",
"secondhand"
],
"shop/sewing":[
"symaskin",
"tyg",
"sy",
"garn",
"Sybutik",
"nå",
"sybutik. sömnadsbutik",
"tråd",
"sömnad"
],
"shop/shoes":[
"Skoaffär",
"skobutik",
"skor"
],
"shop/sports":[
"sportutrustning",
"träningsutrustning",
"träningskläder",
"sportkläder",
"löpskor",
"Sportaffär",
"träningsskor"
],
"shop/stationery":[
"Kontorsmaterial",
"grattiskort",
"papper",
"kort",
"kuvert",
"pennor",
"anteckningsböcker",
"pappersvaror",
"pappershandel",
"Pappershandel"
],
"shop/storage_rental":[
"förråd",
"långtidslager",
"förrådsutrymme",
"bilförvaring",
"magasinera",
"Magasinering",
"förvaring",
"husvagnsförvaring",
"Hyrlager",
"båtförvaring",
"säsongsförvaring",
"vinterförvaring",
"möbelförvaring"
],
"shop/supermarket":[
"supermarket",
"mat",
"snabbköp",
"självbetjäningsbutik",
"Snabbköp",
"affär",
"livsmedelsbutik",
"mataffär",
"självköp",
"dagligvarubutik",
"livsmedel"
],
"shop/tailor":[
"kostym",
"klänning",
"Skräddare",
"kläder"
],
"shop/tattoo":[
"Tatueringsstudio",
"tatuera",
"tatuering",
"tatueringssalong",
"tatuerare"
],
"shop/tea":[
"the",
"Te",
"te",
"teblad",
"thé",
"örtte",
"Te-butik",
"påste"
],
"shop/ticket":[
"biljettlucka",
"biljettkassa",
"biljettkontor",
"Biljettförsäljning",
"biljetter",
"biljettsäljare",
"biljettåterförsäljare"
],
"shop/tiles":[
"kakelplatta",
"plattsättare",
"Klinker",
"plattor",
"Kakelbutik",
"kakel"
],
"shop/tobacco":[
"pipor",
"cigarett",
"röktillbehör",
"tobak",
"cigarr",
"Tobaksbutik",
"cigaretter",
"snus",
"rökning",
"pipa",
"cigarrer"
],
"shop/toys":[
"leksaker",
"barnsaker",
"Leksaksaffär"
],
"shop/trade":[
"Proffshandel",
"granngården",
"trävaror",
"fönster",
"kakel",
"jordbruksprodukter",
"proffsmarknad",
"VVS",
"Trähandel",
"jordbruk",
"brädor",
"byggmaterial",
"lantmannaföreningen",
"brädgård",
"VVS-specialist",
"byggnadsmaterial",
"proffs"
],
"shop/travel_agency":[
"charterflyg",
"charter",
"reseagent",
"Resebyrå",
"biljettförsäljning",
"charterresa"
],
"shop/tyres":[
"däckförsäljning",
"däckbyte",
"hjulbyte",
"fälgar",
"däck",
"fälg",
"hjul",
"Däckfirma",
"hjulförsäljning",
"balansering"
],
"shop/vacant":[
"Tom lokal"
],
"shop/vacuum_cleaner":[
"dammsugaråterförsäljare",
"dammsugarpåsar",
"Dammsugarbutik",
"dammsugartillbehör",
"dammsugare"
],
"shop/variety_store":[
"Fyndbutik",
"överskott",
"lågprisbutik",
"fynd",
"billigt",
"lågpris",
"överskottsaffär"
],
"shop/video":[
"VHS",
"filmbutik",
"filmförsäljning",
"DVD",
"Videobutik",
"filmuthyrning"
],
"shop/video_games":[
"tvspel",
"TV-spel",
"konsolspel",
"spelkonsoler",
"datorspel",
"videospel",
"dataspel"
],
"shop/watches":[
"Klockaffär",
"klockbutik",
"klocka",
"klockor",
"uraffär",
"urbutik",
"ur"
],
"shop/water_sports":[
"Vattensport",
"simning",
"badkläder",
"Vattensport/simning "
],
"shop/weapons":[
"ammunition",
"jakt",
"skjutvapen",
"vapen",
"kniv",
"knivar",
"pistol",
"Vapenaffär"
],
"shop/wholesale":[
"grosshandel",
"grossistverksamhet",
"engros",
"mängdhandel",
"Partihandel",
"lagerklubb",
"grosist",
"Grosistaffär",
"grossistklubb",
"grossistlager"
],
"shop/window_blind":[
"spjälgardin",
"spjäljalusi",
"Persienner",
"markis",
"jalusi",
"rullgardin"
],
"shop/wine":[
"systemet",
"systembolaget",
"vin",
"Vinaffär",
"vinförsäljning"
],
"tourism":[
"turistmagnat",
"turistattraktion",
"Turism",
"sevärdhet"
],
"tourism/alpine_hut":[
"Fjällstuga",
"Fjällstation",
"fjällstation"
],
"tourism/apartment":[
"turist",
"hotell",
"Andelslägenhet",
"Gästlägenhet",
"Turistlägenhet",
"condo",
"lägenhetshotell",
"lägenhet"
],
"tourism/aquarium":[
"fisk",
"Akvarium",
"hav",
"vatten"
],
"tourism/artwork":[
"Publik konst",
"målning",
"gatukonst",
"väggmålning",
"Konst",
"offentlig konst",
"publik konst",
"skulptur",
"staty"
],
"tourism/artwork/mural":[
"fresco",
"mural",
"målning",
"Väggmålning",
"väggmålning"
],
"tourism/artwork/sculpture":[
"Staty",
"byst",
"Skulptur",
"monument",
"snideri",
"skulptur",
"figur"
],
"tourism/artwork/statue":[
"Staty",
"byst",
"monument",
"snideri",
"skulptur",
"figur"
],
"tourism/attraction":[
"Turistattraktion",
"sevärdighet",
"sevärdhet"
],
"tourism/camp_site":[
"tält",
"campinganläggning",
"camping",
"husvagn",
"Campingplats"
],
"tourism/caravan_site":[
"camping",
"husvagnscamping",
"husbilscamping",
"Ställplats",
"campingplats",
"fricamping"
],
"tourism/chalet":[
"helgboende",
"camping",
"stuga",
"sommarstuga",
"Stuga",
"helg",
"semester",
"semesterboende",
"semesterstuga",
"ledighet",
"Campingstuga"
],
"tourism/gallery":[
"Konstgalleri",
"konstverk",
"Konstaffär",
"tavlor",
"kulturer",
"konst",
"konsthandlare",
"konstgalleri",
"galleri",
"statyer",
"konstutställning"
],
"tourism/guest_house":[
"B&D",
"vandrarhem",
"logi",
"övernattningsställe",
"pensionat",
"Bed & Breakfast",
"Gästhus"
],
"tourism/hostel":[
"Vandrarhem",
"övernattningsställe"
],
"tourism/hotel":[
"värdshus",
"Hotell",
"hotellanläggning"
],
"tourism/information":[
"infokarta",
"karta",
"informationskarta",
"Informationstavla",
"Turistbyråer",
"Information",
"turistkontor",
"informationskällan"
],
"tourism/information/board":[
"turistinformation",
"avgång*",
"kollektivtrafik",
"fakta",
"karta",
"Informationstavla",
"information",
"historisk information"
],
"tourism/information/guidepost":[
"Vägmärke",
"Guidepost",
"stigvisning",
"Vägvisare",
"vandringsskyllt"
],
"tourism/information/map":[
"*karta",
"cykelkarta",
"Karta",
"navigering",
"information",
"stadskarta",
"vägkarta",
"informationstavla",
"industrikarta"
],
"tourism/information/office":[
"Turistbyrå",
"turist",
"turistinformation",
"resebyrå",
"turism",
"turistkontor"
],
"tourism/motel":[
"motorhotell",
"hotell",
"väghotell",
"Motell",
"Motel"
],
"tourism/museum":[
"samling",
"museibyggnad",
"historia",
"museum",
"vetenskap",
"utställning",
"konstsamling",
"Museum",
"historik",
"konst",
"arkeologi",
"galleri"
],
"tourism/picnic_site":[
"Picknickplats",
"camping",
"rastplats",
"utflykt",
"campingplats",
"picknick"
],
"tourism/theme_park":[
"nöjespark",
"åkattraktioner",
"nöjesplats",
"tivoli",
"nöjesfält",
"Nöjespark",
"Temapark"
],
"tourism/trail_riding_station":[
"tur",
"ridstation",
"hästrastning",
"häststall",
"gästhus",
"ridningsstation",
"stall",
"turridning",
"Turridningsstation",
"häst"
],
"tourism/viewpoint":[
"utsikt",
"vy",
"Utsiktspunkt",
"Utsiktsplats"
],
"tourism/wilderness_hut":[
"hydda",
"vandring",
"stuga",
"skydd",
"koja",
"hajk",
"kyffe",
"övernattning",
"Stuga (för vandrare o.d.)",
"vildmarksstuga",
"barack",
"fjällstuga",
"fjällstation",
"Ödestuga"
],
"tourism/zoo":[
"djurpark",
"Zoo",
"zoologisk trädgård"
],
"traffic_calming":[
"långsam",
"hastighet",
"fartgupp",
"* fart*",
"gupp",
"trafikhinder",
"säkerhet",
"Farthinder"
],
"traffic_calming/bump":[
"bula",
"Fartbula (kort gupp)",
"bump",
"fartgupp",
"vägbula",
"farthinder",
"Fartbula",
"gupp"
],
"traffic_calming/chicane":[
"trafikchikan",
"långsam",
"hastighet",
"* fart*",
"Sidoförskjutning (chikan)",
"kurvor",
"Sidoförskjutning",
"chikan",
"slalom",
"trafikhinder",
"säkerhet",
"Farthinder"
],
"traffic_calming/choker":[
"lins",
"choker",
"Avsmalning",
"Timglas",
"långsam",
"hastighet",
"* fart*",
"trafikhinder",
"Farthinder",
"säkerhet"
],
"traffic_calming/cushion":[
"Timglas",
"långsam",
"hastighet",
"Vägkudde",
"Farthinder",
"lins",
"vägkudde",
"fartgupp",
"* fart*",
"farthinder",
"trafikhinder",
"gupp",
"säkerhet"
],
"traffic_calming/dip":[
"långsam",
"hastighet",
"fartgupp",
"grop",
"* fart*",
"farthinder",
"trafikhinder",
"Grop",
"Farthinder",
"säkerhet",
"försänkning"
],
"traffic_calming/hump":[
"Wattgupp",
"normalt fartgupp",
"Wattska guppet",
"fartpuckel",
"GP-gupp",
"puckel",
"fartgupp",
"farthinder",
"Normalt fartgupp",
"Cirkulärt gupp",
"standardgupp",
"gupp"
],
"traffic_calming/island":[
"cirkulation",
"långsam",
"hastighet",
"cirkel",
"sidorefug",
"Farthinder",
"mittrefug",
"trafikö",
"ö",
"Refug",
"cirkulationsplats",
"* fart*",
"farthinder",
"trafikhinder",
"säkerhet",
"rondell"
],
"traffic_calming/rumble_strip":[
"Bullerräfflor",
"Pennsylvaniaräfflor"
],
"traffic_calming/table":[
"Fartgupp (långt)",
"fartgupp",
"farthinder",
"långt fartgupp",
"gupp",
"Platågupp"
],
"traffic_sign":[
"Trafikskyllt",
"Vägmärke",
"trafikmärke",
"skyllt",
"vägskyllt",
"vägmärke",
"vägvisare"
],
"traffic_sign/city_limit":[
"Skyllt för tättbebyggt område",
"skyllt",
"Tättbebyggt område",
"stadsgräns",
"ort",
"Trafikskyllt",
"stad",
"tätort",
"trafikmärke",
"gräns",
"vägskyllt",
"vägmärke",
"vägvisare"
],
"traffic_sign/city_limit_vertex":[
"Skyllt för tättbebyggt område",
"skyllt",
"Tättbebyggt område",
"stadsgräns",
"ort",
"Trafikskyllt",
"stad",
"tätort",
"trafikmärke",
"gräns",
"vägskyllt",
"vägmärke",
"vägvisare"
],
"traffic_sign/maxspeed":[
"Trafikskyllt",
"fart",
"maxhastighet",
"trafikmärke",
"maxfart",
"skyllt",
"hastighet",
"Hastighetsskylt",
"Hastighetsbegränsning",
"vägskyllt",
"vägmärke",
"vägvisare"
],
"traffic_sign/maxspeed_vertex":[
"Trafikskyllt",
"fart",
"maxhastighet",
"trafikmärke",
"maxfart",
"skyllt",
"hastighet",
"Hastighetsskylt",
"Hastighetsbegränsning",
"vägskyllt",
"vägmärke",
"vägvisare"
],
"traffic_sign_vertex":[
"Trafikskyllt",
"Vägmärke",
"trafikmärke",
"skyllt",
"vägskyllt",
"vägmärke",
"vägvisare"
],
"type/boundary":[
"Gräns",
"gränslinje",
"administrativ gräns"
],
"type/boundary/administrative":[
"Administrativ gräns",
"stat",
"administrativ enhet",
"gräns",
"territorium"
],
"type/multipolygon":[
"Multipolygon"
],
"type/restriction":[
"begränsning",
"inskränkning",
"Restriktion",
"förbehåll"
],
"type/restriction/no_left_turn":[
"Ingen vänstersväng",
"sväng ej vänster"
],
"type/restriction/no_right_turn":[
"ej högersväng",
"Ingen högersväng",
"sväng ej höger"
],
"type/restriction/no_straight_on":[
"ej rakt fram",
"Ej rakt fram",
"Fortsätt ej framåt"
],
"type/restriction/no_u_turn":[
"får ej vända",
"Ingen U-sväng"
],
"type/restriction/only_left_turn":[
"vänster",
"Enbart vänstersväng",
"vänstersväng"
],
"type/restriction/only_right_turn":[
"Enbart högersväng",
"högersväng",
"höger"
],
"type/restriction/only_straight_on":[
"Enbart rakt fram",
"fortsätt framåt",
"får ej svänga"
],
"type/restriction/only_u_turn":[
"måste vända",
"U-sväng",
"Enbart U-sväng"
],
"type/route":[
"Rutt",
"rutt",
"färdled",
"färdväg"
],
"type/route/bicycle":[
"cykelled",
"cykelförbindelse",
"cykelnät",
"Cykelrutt"
],
"type/route/bus":[
"busslinje",
"bussväg",
"Busslinje",
"Bussrutt",
"bussled"
],
"type/route/detour":[
"Alternativ rutt",
"omväg",
"alternativ väg"
],
"type/route/ferry":[
"båtrutt",
"båtlinjetrafik",
"Färjerutt"
],
"type/route/foot":[
"Vandringsled",
"vandringsled",
"stig",
"Vandringsrutt"
],
"type/route/hiking":[
"Vandringsled",
"vandringsled",
"stig",
"Vandringsrutt"
],
"type/route/horse":[
"Hästspår",
"rida",
"Ridrutt",
"ridning",
"hästspår",
"hästrutt",
"ridspår",
"häst"
],
"type/route/light_rail":[
"tågrutt",
"smalspårig järnväg",
"rutt för snabbspårväg",
"järnvägsförbindelse",
"stadsbana",
"järnvägsrutt",
"snabbspårväg",
"smalspår",
"Rutt på snabbspårväg / stadsbana",
"tågnät",
"rutt för stadsbana",
"Rutt på smalspårig järnväg",
"järnväg"
],
"type/route/pipeline":[
"pipeline",
"oljeledning",
"vattenledning",
"avloppsledning",
"rörledning",
"Rörledningsrutt"
],
"type/route/piste":[
"längdskidspår",
"pistspår",
"Pist/skidrutt",
"skidor",
"skidtur",
"snöpark",
"skidbacke",
"utförsåkning",
"skridskorutt",
"skidrutt",
"slädspår",
"längdskidåkning",
"slalombacke",
"skidspår",
"skidbana",
"skridskospår",
"skridskobana",
"Pist"
],
"type/route/power":[
"kraftledning",
"elnät",
"Kraftledningsrutt",
"elförsörjning"
],
"type/route/road":[
"Vägrutt",
"vägförbindelse",
"vägnät"
],
"type/route/subway":[
"Tunnelbanerutt",
"tunnelbana"
],
"type/route/train":[
"tågnät",
"järnvägsförbindelse",
"Tågrutt",
"järnväg",
"järnvägsrutt"
],
"type/route/tram":[
"spårvagnsnät",
"Spårvagnsrutt",
"spårvagn",
"spårvagnsförbindelse",
"spårvagnsräls"
],
"type/route_master":[
"huvudförbindelse",
"Huvudrutt",
"huvudväg"
],
"type/site":[
"anläggning",
"läge",
"ställe",
"Plats"
],
"type/waterway":[
"Vattenväg",
"vattendrag",
"Vattendrag",
"vattenflöde"
],
"vertex":[
"Annat",
"övrigt"
],
"waterway":[
"Vattenväg"
],
"waterway/boatyard":[
"båtställplats",
"varv",
"Båtvarv",
"uppläggningsplats",
"vinterförvaring"
],
"waterway/canal":[
"vattenväg",
"vattenled",
"Kanal"
],
"waterway/dam":[
"fördämning",
"vattensamling",
"damm",
"reservoar",
"Fördämning"
],
"waterway/ditch":[
"Dike",
"fåra"
],
"waterway/dock":[
"båtdocka",
"båtvarv",
"fartygsvarv",
"Våt- / Torrdocka",
"varv",
"Torrdocka",
"docka",
"lastdocka",
"våtdocka",
"fartygsdocka"
],
"waterway/drain":[
"dagvattenavrinning",
"dagvatten",
"Dränering",
"dränering",
"avrinning"
],
"waterway/fuel":[
"båtmack",
"tankstation båtbensninmack",
"bränslestation",
"båtmensinstation",
"Sjömack"
],
"waterway/milestone":[
"Milsten vid vattendrag",
"kilometertavla",
"kilometerpåle",
"sjöfart",
"milsten",
"referenstavla",
"kilometerstolpe",
"avståndsmärke"
],
"waterway/river":[
"vattendrag",
"ström",
"jokk",
"Å",
"fors",
"Flod",
"flod",
"älv"
],
"waterway/riverbank":[
"åstrand",
"flodbank",
"flodstrand",
"Flodbank"
],
"waterway/sanitary_dump_station":[
"tömningsplats",
"båtlatrin",
"CTDP",
"Dumpstation",
"gråvatten",
"båtsanitet",
"gråvattentömning",
"Elsan",
"Marin latrintömning",
"sanitet",
"Pumpa ut",
"latrintömning",
"CDP",
"båttömnig",
"Båt",
"sanitära",
"kemisk toalett",
"toalettömning",
"utpumpning",
"campingtoalett",
"Vattenfarkoster"
],
"waterway/stream":[
"dike",
"biflod",
"vattendrag",
"flöde",
"ström",
"bäck",
"biflöde",
"flod",
"Bäck",
"rännil"
],
"waterway/stream_intermittent":[
"Arroyo",
"Periodiskt vattendrag",
"bäck",
"periodiskt",
"dagvatten",
"biflöde",
"tillfälligt",
"översvämning",
"dike",
"vattendrag",
"tillfälligt vattendrag",
"dränering",
"avrinning",
"rännil"
],
"waterway/water_point":[
"Dricksvatten",
"Dricksvatten för båt",
"vattenpåfyllning",
"vattentank"
],
"waterway/waterfall":[
"Vattenfall",
"fall",
"fors"
],
"waterway/weir":[
"fördämning",
"vattensamling",
"damm",
"reservoar",
"Damm"
]
}
